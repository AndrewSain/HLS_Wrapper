
// Register/Wire Declarations

reg [5:0] reg_time_i[0:6][0:8][0:1];
reg [1:0] reg_vl_i[0:12][0:8];
reg [3:0] reg_q_i[0:12][0:8][0:2];
reg [3:0] reg_cpatr_i[0:5][0:8][0:1];
reg [12:0] reg_ph_i[0:5][0:8][0:1];
reg [6:0] reg_th11_i[0:5][0:8][0:1];
reg [6:0] reg_th_i[0:2][0:2][0:3];
reg [6:0] reg_phzvl_i[0:12][0:8];
reg [43:0] reg_ph_hit_i[0:12][0:8];
reg [5:0] reg_time_o[0:0][0:6][0:8][0:1];
reg [1:0] reg_vl_o[0:0][0:12][0:8];
reg [3:0] reg_q_o[0:0][0:12][0:8][0:2];
reg [3:0] reg_cpatr_o[0:0][0:5][0:8][0:1];
reg [12:0] reg_ph_o[0:0][0:5][0:8][0:1];
reg [6:0] reg_th11_o[0:0][0:5][0:8][0:1];
reg [6:0] reg_th_o[0:0][0:2][0:2][0:3];
reg [6:0] reg_phzvl_o[0:0][0:12][0:8];
reg [43:0] reg_ph_hit_o[0:0][0:12][0:8];
wire [5:0] wire_time_o[0:0][0:6][0:8][0:1];
wire [1:0] wire_vl_o[0:0][0:12][0:8];
wire [3:0] wire_q_o[0:0][0:12][0:8][0:2];
wire [3:0] wire_cpatr_o[0:0][0:5][0:8][0:1];
wire [12:0] wire_ph_o[0:0][0:5][0:8][0:1];
wire [6:0] wire_th11_o[0:0][0:5][0:8][0:1];
wire [6:0] wire_th_o[0:0][0:2][0:2][0:3];
wire [6:0] wire_phzvl_o[0:0][0:12][0:8];
wire [43:0] wire_ph_hit_o[0:0][0:12][0:8];

// IO Connections

.time_i_0_0_0_V(reg_time_i[0][0][0]),
.time_i_0_0_1_V(reg_time_i[0][0][1]),
.time_i_0_1_0_V(reg_time_i[0][1][0]),
.time_i_0_1_1_V(reg_time_i[0][1][1]),
.time_i_0_2_0_V(reg_time_i[0][2][0]),
.time_i_0_2_1_V(reg_time_i[0][2][1]),
.time_i_0_3_0_V(reg_time_i[0][3][0]),
.time_i_0_3_1_V(reg_time_i[0][3][1]),
.time_i_0_4_0_V(reg_time_i[0][4][0]),
.time_i_0_4_1_V(reg_time_i[0][4][1]),
.time_i_0_5_0_V(reg_time_i[0][5][0]),
.time_i_0_5_1_V(reg_time_i[0][5][1]),
.time_i_0_6_0_V(reg_time_i[0][6][0]),
.time_i_0_6_1_V(reg_time_i[0][6][1]),
.time_i_0_7_0_V(reg_time_i[0][7][0]),
.time_i_0_7_1_V(reg_time_i[0][7][1]),
.time_i_0_8_0_V(reg_time_i[0][8][0]),
.time_i_0_8_1_V(reg_time_i[0][8][1]),
.time_i_1_0_0_V(reg_time_i[1][0][0]),
.time_i_1_0_1_V(reg_time_i[1][0][1]),
.time_i_1_1_0_V(reg_time_i[1][1][0]),
.time_i_1_1_1_V(reg_time_i[1][1][1]),
.time_i_1_2_0_V(reg_time_i[1][2][0]),
.time_i_1_2_1_V(reg_time_i[1][2][1]),
.time_i_1_3_0_V(reg_time_i[1][3][0]),
.time_i_1_3_1_V(reg_time_i[1][3][1]),
.time_i_1_4_0_V(reg_time_i[1][4][0]),
.time_i_1_4_1_V(reg_time_i[1][4][1]),
.time_i_1_5_0_V(reg_time_i[1][5][0]),
.time_i_1_5_1_V(reg_time_i[1][5][1]),
.time_i_1_6_0_V(reg_time_i[1][6][0]),
.time_i_1_6_1_V(reg_time_i[1][6][1]),
.time_i_1_7_0_V(reg_time_i[1][7][0]),
.time_i_1_7_1_V(reg_time_i[1][7][1]),
.time_i_1_8_0_V(reg_time_i[1][8][0]),
.time_i_1_8_1_V(reg_time_i[1][8][1]),
.time_i_2_0_0_V(reg_time_i[2][0][0]),
.time_i_2_0_1_V(reg_time_i[2][0][1]),
.time_i_2_1_0_V(reg_time_i[2][1][0]),
.time_i_2_1_1_V(reg_time_i[2][1][1]),
.time_i_2_2_0_V(reg_time_i[2][2][0]),
.time_i_2_2_1_V(reg_time_i[2][2][1]),
.time_i_2_3_0_V(reg_time_i[2][3][0]),
.time_i_2_3_1_V(reg_time_i[2][3][1]),
.time_i_2_4_0_V(reg_time_i[2][4][0]),
.time_i_2_4_1_V(reg_time_i[2][4][1]),
.time_i_2_5_0_V(reg_time_i[2][5][0]),
.time_i_2_5_1_V(reg_time_i[2][5][1]),
.time_i_2_6_0_V(reg_time_i[2][6][0]),
.time_i_2_6_1_V(reg_time_i[2][6][1]),
.time_i_2_7_0_V(reg_time_i[2][7][0]),
.time_i_2_7_1_V(reg_time_i[2][7][1]),
.time_i_2_8_0_V(reg_time_i[2][8][0]),
.time_i_2_8_1_V(reg_time_i[2][8][1]),
.time_i_3_0_0_V(reg_time_i[3][0][0]),
.time_i_3_0_1_V(reg_time_i[3][0][1]),
.time_i_3_1_0_V(reg_time_i[3][1][0]),
.time_i_3_1_1_V(reg_time_i[3][1][1]),
.time_i_3_2_0_V(reg_time_i[3][2][0]),
.time_i_3_2_1_V(reg_time_i[3][2][1]),
.time_i_3_3_0_V(reg_time_i[3][3][0]),
.time_i_3_3_1_V(reg_time_i[3][3][1]),
.time_i_3_4_0_V(reg_time_i[3][4][0]),
.time_i_3_4_1_V(reg_time_i[3][4][1]),
.time_i_3_5_0_V(reg_time_i[3][5][0]),
.time_i_3_5_1_V(reg_time_i[3][5][1]),
.time_i_3_6_0_V(reg_time_i[3][6][0]),
.time_i_3_6_1_V(reg_time_i[3][6][1]),
.time_i_3_7_0_V(reg_time_i[3][7][0]),
.time_i_3_7_1_V(reg_time_i[3][7][1]),
.time_i_3_8_0_V(reg_time_i[3][8][0]),
.time_i_3_8_1_V(reg_time_i[3][8][1]),
.time_i_4_0_0_V(reg_time_i[4][0][0]),
.time_i_4_0_1_V(reg_time_i[4][0][1]),
.time_i_4_1_0_V(reg_time_i[4][1][0]),
.time_i_4_1_1_V(reg_time_i[4][1][1]),
.time_i_4_2_0_V(reg_time_i[4][2][0]),
.time_i_4_2_1_V(reg_time_i[4][2][1]),
.time_i_4_3_0_V(reg_time_i[4][3][0]),
.time_i_4_3_1_V(reg_time_i[4][3][1]),
.time_i_4_4_0_V(reg_time_i[4][4][0]),
.time_i_4_4_1_V(reg_time_i[4][4][1]),
.time_i_4_5_0_V(reg_time_i[4][5][0]),
.time_i_4_5_1_V(reg_time_i[4][5][1]),
.time_i_4_6_0_V(reg_time_i[4][6][0]),
.time_i_4_6_1_V(reg_time_i[4][6][1]),
.time_i_4_7_0_V(reg_time_i[4][7][0]),
.time_i_4_7_1_V(reg_time_i[4][7][1]),
.time_i_4_8_0_V(reg_time_i[4][8][0]),
.time_i_4_8_1_V(reg_time_i[4][8][1]),
.time_i_5_0_0_V(reg_time_i[5][0][0]),
.time_i_5_0_1_V(reg_time_i[5][0][1]),
.time_i_5_1_0_V(reg_time_i[5][1][0]),
.time_i_5_1_1_V(reg_time_i[5][1][1]),
.time_i_5_2_0_V(reg_time_i[5][2][0]),
.time_i_5_2_1_V(reg_time_i[5][2][1]),
.time_i_5_3_0_V(reg_time_i[5][3][0]),
.time_i_5_3_1_V(reg_time_i[5][3][1]),
.time_i_5_4_0_V(reg_time_i[5][4][0]),
.time_i_5_4_1_V(reg_time_i[5][4][1]),
.time_i_5_5_0_V(reg_time_i[5][5][0]),
.time_i_5_5_1_V(reg_time_i[5][5][1]),
.time_i_5_6_0_V(reg_time_i[5][6][0]),
.time_i_5_6_1_V(reg_time_i[5][6][1]),
.time_i_5_7_0_V(reg_time_i[5][7][0]),
.time_i_5_7_1_V(reg_time_i[5][7][1]),
.time_i_5_8_0_V(reg_time_i[5][8][0]),
.time_i_5_8_1_V(reg_time_i[5][8][1]),
.time_i_6_0_0_V(reg_time_i[6][0][0]),
.time_i_6_0_1_V(reg_time_i[6][0][1]),
.time_i_6_1_0_V(reg_time_i[6][1][0]),
.time_i_6_1_1_V(reg_time_i[6][1][1]),
.time_i_6_2_0_V(reg_time_i[6][2][0]),
.time_i_6_2_1_V(reg_time_i[6][2][1]),
.time_i_6_3_0_V(reg_time_i[6][3][0]),
.time_i_6_3_1_V(reg_time_i[6][3][1]),
.time_i_6_4_0_V(reg_time_i[6][4][0]),
.time_i_6_4_1_V(reg_time_i[6][4][1]),
.time_i_6_5_0_V(reg_time_i[6][5][0]),
.time_i_6_5_1_V(reg_time_i[6][5][1]),
.time_i_6_6_0_V(reg_time_i[6][6][0]),
.time_i_6_6_1_V(reg_time_i[6][6][1]),
.time_i_6_7_0_V(reg_time_i[6][7][0]),
.time_i_6_7_1_V(reg_time_i[6][7][1]),
.time_i_6_8_0_V(reg_time_i[6][8][0]),
.time_i_6_8_1_V(reg_time_i[6][8][1]),
.vl_i_0_0_V(reg_vl_i[0][0]),
.vl_i_0_1_V(reg_vl_i[0][1]),
.vl_i_0_2_V(reg_vl_i[0][2]),
.vl_i_0_3_V(reg_vl_i[0][3]),
.vl_i_0_4_V(reg_vl_i[0][4]),
.vl_i_0_5_V(reg_vl_i[0][5]),
.vl_i_0_6_V(reg_vl_i[0][6]),
.vl_i_0_7_V(reg_vl_i[0][7]),
.vl_i_0_8_V(reg_vl_i[0][8]),
.vl_i_1_0_V(reg_vl_i[1][0]),
.vl_i_1_1_V(reg_vl_i[1][1]),
.vl_i_1_2_V(reg_vl_i[1][2]),
.vl_i_1_3_V(reg_vl_i[1][3]),
.vl_i_1_4_V(reg_vl_i[1][4]),
.vl_i_1_5_V(reg_vl_i[1][5]),
.vl_i_1_6_V(reg_vl_i[1][6]),
.vl_i_1_7_V(reg_vl_i[1][7]),
.vl_i_1_8_V(reg_vl_i[1][8]),
.vl_i_2_0_V(reg_vl_i[2][0]),
.vl_i_2_1_V(reg_vl_i[2][1]),
.vl_i_2_2_V(reg_vl_i[2][2]),
.vl_i_2_3_V(reg_vl_i[2][3]),
.vl_i_2_4_V(reg_vl_i[2][4]),
.vl_i_2_5_V(reg_vl_i[2][5]),
.vl_i_2_6_V(reg_vl_i[2][6]),
.vl_i_2_7_V(reg_vl_i[2][7]),
.vl_i_2_8_V(reg_vl_i[2][8]),
.vl_i_3_0_V(reg_vl_i[3][0]),
.vl_i_3_1_V(reg_vl_i[3][1]),
.vl_i_3_2_V(reg_vl_i[3][2]),
.vl_i_3_3_V(reg_vl_i[3][3]),
.vl_i_3_4_V(reg_vl_i[3][4]),
.vl_i_3_5_V(reg_vl_i[3][5]),
.vl_i_3_6_V(reg_vl_i[3][6]),
.vl_i_3_7_V(reg_vl_i[3][7]),
.vl_i_3_8_V(reg_vl_i[3][8]),
.vl_i_4_0_V(reg_vl_i[4][0]),
.vl_i_4_1_V(reg_vl_i[4][1]),
.vl_i_4_2_V(reg_vl_i[4][2]),
.vl_i_4_3_V(reg_vl_i[4][3]),
.vl_i_4_4_V(reg_vl_i[4][4]),
.vl_i_4_5_V(reg_vl_i[4][5]),
.vl_i_4_6_V(reg_vl_i[4][6]),
.vl_i_4_7_V(reg_vl_i[4][7]),
.vl_i_4_8_V(reg_vl_i[4][8]),
.vl_i_5_0_V(reg_vl_i[5][0]),
.vl_i_5_1_V(reg_vl_i[5][1]),
.vl_i_5_2_V(reg_vl_i[5][2]),
.vl_i_5_3_V(reg_vl_i[5][3]),
.vl_i_5_4_V(reg_vl_i[5][4]),
.vl_i_5_5_V(reg_vl_i[5][5]),
.vl_i_5_6_V(reg_vl_i[5][6]),
.vl_i_5_7_V(reg_vl_i[5][7]),
.vl_i_5_8_V(reg_vl_i[5][8]),
.vl_i_6_0_V(reg_vl_i[6][0]),
.vl_i_6_1_V(reg_vl_i[6][1]),
.vl_i_6_2_V(reg_vl_i[6][2]),
.vl_i_6_3_V(reg_vl_i[6][3]),
.vl_i_6_4_V(reg_vl_i[6][4]),
.vl_i_6_5_V(reg_vl_i[6][5]),
.vl_i_6_6_V(reg_vl_i[6][6]),
.vl_i_6_7_V(reg_vl_i[6][7]),
.vl_i_6_8_V(reg_vl_i[6][8]),
.vl_i_7_0_V(reg_vl_i[7][0]),
.vl_i_7_1_V(reg_vl_i[7][1]),
.vl_i_7_2_V(reg_vl_i[7][2]),
.vl_i_7_3_V(reg_vl_i[7][3]),
.vl_i_7_4_V(reg_vl_i[7][4]),
.vl_i_7_5_V(reg_vl_i[7][5]),
.vl_i_7_6_V(reg_vl_i[7][6]),
.vl_i_7_7_V(reg_vl_i[7][7]),
.vl_i_7_8_V(reg_vl_i[7][8]),
.vl_i_8_0_V(reg_vl_i[8][0]),
.vl_i_8_1_V(reg_vl_i[8][1]),
.vl_i_8_2_V(reg_vl_i[8][2]),
.vl_i_8_3_V(reg_vl_i[8][3]),
.vl_i_8_4_V(reg_vl_i[8][4]),
.vl_i_8_5_V(reg_vl_i[8][5]),
.vl_i_8_6_V(reg_vl_i[8][6]),
.vl_i_8_7_V(reg_vl_i[8][7]),
.vl_i_8_8_V(reg_vl_i[8][8]),
.vl_i_9_0_V(reg_vl_i[9][0]),
.vl_i_9_1_V(reg_vl_i[9][1]),
.vl_i_9_2_V(reg_vl_i[9][2]),
.vl_i_9_3_V(reg_vl_i[9][3]),
.vl_i_9_4_V(reg_vl_i[9][4]),
.vl_i_9_5_V(reg_vl_i[9][5]),
.vl_i_9_6_V(reg_vl_i[9][6]),
.vl_i_9_7_V(reg_vl_i[9][7]),
.vl_i_9_8_V(reg_vl_i[9][8]),
.vl_i_10_0_V(reg_vl_i[10][0]),
.vl_i_10_1_V(reg_vl_i[10][1]),
.vl_i_10_2_V(reg_vl_i[10][2]),
.vl_i_10_3_V(reg_vl_i[10][3]),
.vl_i_10_4_V(reg_vl_i[10][4]),
.vl_i_10_5_V(reg_vl_i[10][5]),
.vl_i_10_6_V(reg_vl_i[10][6]),
.vl_i_10_7_V(reg_vl_i[10][7]),
.vl_i_10_8_V(reg_vl_i[10][8]),
.vl_i_11_0_V(reg_vl_i[11][0]),
.vl_i_11_1_V(reg_vl_i[11][1]),
.vl_i_11_2_V(reg_vl_i[11][2]),
.vl_i_11_3_V(reg_vl_i[11][3]),
.vl_i_11_4_V(reg_vl_i[11][4]),
.vl_i_11_5_V(reg_vl_i[11][5]),
.vl_i_11_6_V(reg_vl_i[11][6]),
.vl_i_11_7_V(reg_vl_i[11][7]),
.vl_i_11_8_V(reg_vl_i[11][8]),
.vl_i_12_0_V(reg_vl_i[12][0]),
.vl_i_12_1_V(reg_vl_i[12][1]),
.vl_i_12_2_V(reg_vl_i[12][2]),
.vl_i_12_3_V(reg_vl_i[12][3]),
.vl_i_12_4_V(reg_vl_i[12][4]),
.vl_i_12_5_V(reg_vl_i[12][5]),
.vl_i_12_6_V(reg_vl_i[12][6]),
.vl_i_12_7_V(reg_vl_i[12][7]),
.vl_i_12_8_V(reg_vl_i[12][8]),
.q_i_0_0_0_V(reg_q_i[0][0][0]),
.q_i_0_0_1_V(reg_q_i[0][0][1]),
.q_i_0_0_2_V(reg_q_i[0][0][2]),
.q_i_0_1_0_V(reg_q_i[0][1][0]),
.q_i_0_1_1_V(reg_q_i[0][1][1]),
.q_i_0_1_2_V(reg_q_i[0][1][2]),
.q_i_0_2_0_V(reg_q_i[0][2][0]),
.q_i_0_2_1_V(reg_q_i[0][2][1]),
.q_i_0_2_2_V(reg_q_i[0][2][2]),
.q_i_0_3_0_V(reg_q_i[0][3][0]),
.q_i_0_3_1_V(reg_q_i[0][3][1]),
.q_i_0_3_2_V(reg_q_i[0][3][2]),
.q_i_0_4_0_V(reg_q_i[0][4][0]),
.q_i_0_4_1_V(reg_q_i[0][4][1]),
.q_i_0_4_2_V(reg_q_i[0][4][2]),
.q_i_0_5_0_V(reg_q_i[0][5][0]),
.q_i_0_5_1_V(reg_q_i[0][5][1]),
.q_i_0_5_2_V(reg_q_i[0][5][2]),
.q_i_0_6_0_V(reg_q_i[0][6][0]),
.q_i_0_6_1_V(reg_q_i[0][6][1]),
.q_i_0_6_2_V(reg_q_i[0][6][2]),
.q_i_0_7_0_V(reg_q_i[0][7][0]),
.q_i_0_7_1_V(reg_q_i[0][7][1]),
.q_i_0_7_2_V(reg_q_i[0][7][2]),
.q_i_0_8_0_V(reg_q_i[0][8][0]),
.q_i_0_8_1_V(reg_q_i[0][8][1]),
.q_i_0_8_2_V(reg_q_i[0][8][2]),
.q_i_1_0_0_V(reg_q_i[1][0][0]),
.q_i_1_0_1_V(reg_q_i[1][0][1]),
.q_i_1_0_2_V(reg_q_i[1][0][2]),
.q_i_1_1_0_V(reg_q_i[1][1][0]),
.q_i_1_1_1_V(reg_q_i[1][1][1]),
.q_i_1_1_2_V(reg_q_i[1][1][2]),
.q_i_1_2_0_V(reg_q_i[1][2][0]),
.q_i_1_2_1_V(reg_q_i[1][2][1]),
.q_i_1_2_2_V(reg_q_i[1][2][2]),
.q_i_1_3_0_V(reg_q_i[1][3][0]),
.q_i_1_3_1_V(reg_q_i[1][3][1]),
.q_i_1_3_2_V(reg_q_i[1][3][2]),
.q_i_1_4_0_V(reg_q_i[1][4][0]),
.q_i_1_4_1_V(reg_q_i[1][4][1]),
.q_i_1_4_2_V(reg_q_i[1][4][2]),
.q_i_1_5_0_V(reg_q_i[1][5][0]),
.q_i_1_5_1_V(reg_q_i[1][5][1]),
.q_i_1_5_2_V(reg_q_i[1][5][2]),
.q_i_1_6_0_V(reg_q_i[1][6][0]),
.q_i_1_6_1_V(reg_q_i[1][6][1]),
.q_i_1_6_2_V(reg_q_i[1][6][2]),
.q_i_1_7_0_V(reg_q_i[1][7][0]),
.q_i_1_7_1_V(reg_q_i[1][7][1]),
.q_i_1_7_2_V(reg_q_i[1][7][2]),
.q_i_1_8_0_V(reg_q_i[1][8][0]),
.q_i_1_8_1_V(reg_q_i[1][8][1]),
.q_i_1_8_2_V(reg_q_i[1][8][2]),
.q_i_2_0_0_V(reg_q_i[2][0][0]),
.q_i_2_0_1_V(reg_q_i[2][0][1]),
.q_i_2_0_2_V(reg_q_i[2][0][2]),
.q_i_2_1_0_V(reg_q_i[2][1][0]),
.q_i_2_1_1_V(reg_q_i[2][1][1]),
.q_i_2_1_2_V(reg_q_i[2][1][2]),
.q_i_2_2_0_V(reg_q_i[2][2][0]),
.q_i_2_2_1_V(reg_q_i[2][2][1]),
.q_i_2_2_2_V(reg_q_i[2][2][2]),
.q_i_2_3_0_V(reg_q_i[2][3][0]),
.q_i_2_3_1_V(reg_q_i[2][3][1]),
.q_i_2_3_2_V(reg_q_i[2][3][2]),
.q_i_2_4_0_V(reg_q_i[2][4][0]),
.q_i_2_4_1_V(reg_q_i[2][4][1]),
.q_i_2_4_2_V(reg_q_i[2][4][2]),
.q_i_2_5_0_V(reg_q_i[2][5][0]),
.q_i_2_5_1_V(reg_q_i[2][5][1]),
.q_i_2_5_2_V(reg_q_i[2][5][2]),
.q_i_2_6_0_V(reg_q_i[2][6][0]),
.q_i_2_6_1_V(reg_q_i[2][6][1]),
.q_i_2_6_2_V(reg_q_i[2][6][2]),
.q_i_2_7_0_V(reg_q_i[2][7][0]),
.q_i_2_7_1_V(reg_q_i[2][7][1]),
.q_i_2_7_2_V(reg_q_i[2][7][2]),
.q_i_2_8_0_V(reg_q_i[2][8][0]),
.q_i_2_8_1_V(reg_q_i[2][8][1]),
.q_i_2_8_2_V(reg_q_i[2][8][2]),
.q_i_3_0_0_V(reg_q_i[3][0][0]),
.q_i_3_0_1_V(reg_q_i[3][0][1]),
.q_i_3_0_2_V(reg_q_i[3][0][2]),
.q_i_3_1_0_V(reg_q_i[3][1][0]),
.q_i_3_1_1_V(reg_q_i[3][1][1]),
.q_i_3_1_2_V(reg_q_i[3][1][2]),
.q_i_3_2_0_V(reg_q_i[3][2][0]),
.q_i_3_2_1_V(reg_q_i[3][2][1]),
.q_i_3_2_2_V(reg_q_i[3][2][2]),
.q_i_3_3_0_V(reg_q_i[3][3][0]),
.q_i_3_3_1_V(reg_q_i[3][3][1]),
.q_i_3_3_2_V(reg_q_i[3][3][2]),
.q_i_3_4_0_V(reg_q_i[3][4][0]),
.q_i_3_4_1_V(reg_q_i[3][4][1]),
.q_i_3_4_2_V(reg_q_i[3][4][2]),
.q_i_3_5_0_V(reg_q_i[3][5][0]),
.q_i_3_5_1_V(reg_q_i[3][5][1]),
.q_i_3_5_2_V(reg_q_i[3][5][2]),
.q_i_3_6_0_V(reg_q_i[3][6][0]),
.q_i_3_6_1_V(reg_q_i[3][6][1]),
.q_i_3_6_2_V(reg_q_i[3][6][2]),
.q_i_3_7_0_V(reg_q_i[3][7][0]),
.q_i_3_7_1_V(reg_q_i[3][7][1]),
.q_i_3_7_2_V(reg_q_i[3][7][2]),
.q_i_3_8_0_V(reg_q_i[3][8][0]),
.q_i_3_8_1_V(reg_q_i[3][8][1]),
.q_i_3_8_2_V(reg_q_i[3][8][2]),
.q_i_4_0_0_V(reg_q_i[4][0][0]),
.q_i_4_0_1_V(reg_q_i[4][0][1]),
.q_i_4_0_2_V(reg_q_i[4][0][2]),
.q_i_4_1_0_V(reg_q_i[4][1][0]),
.q_i_4_1_1_V(reg_q_i[4][1][1]),
.q_i_4_1_2_V(reg_q_i[4][1][2]),
.q_i_4_2_0_V(reg_q_i[4][2][0]),
.q_i_4_2_1_V(reg_q_i[4][2][1]),
.q_i_4_2_2_V(reg_q_i[4][2][2]),
.q_i_4_3_0_V(reg_q_i[4][3][0]),
.q_i_4_3_1_V(reg_q_i[4][3][1]),
.q_i_4_3_2_V(reg_q_i[4][3][2]),
.q_i_4_4_0_V(reg_q_i[4][4][0]),
.q_i_4_4_1_V(reg_q_i[4][4][1]),
.q_i_4_4_2_V(reg_q_i[4][4][2]),
.q_i_4_5_0_V(reg_q_i[4][5][0]),
.q_i_4_5_1_V(reg_q_i[4][5][1]),
.q_i_4_5_2_V(reg_q_i[4][5][2]),
.q_i_4_6_0_V(reg_q_i[4][6][0]),
.q_i_4_6_1_V(reg_q_i[4][6][1]),
.q_i_4_6_2_V(reg_q_i[4][6][2]),
.q_i_4_7_0_V(reg_q_i[4][7][0]),
.q_i_4_7_1_V(reg_q_i[4][7][1]),
.q_i_4_7_2_V(reg_q_i[4][7][2]),
.q_i_4_8_0_V(reg_q_i[4][8][0]),
.q_i_4_8_1_V(reg_q_i[4][8][1]),
.q_i_4_8_2_V(reg_q_i[4][8][2]),
.q_i_5_0_0_V(reg_q_i[5][0][0]),
.q_i_5_0_1_V(reg_q_i[5][0][1]),
.q_i_5_0_2_V(reg_q_i[5][0][2]),
.q_i_5_1_0_V(reg_q_i[5][1][0]),
.q_i_5_1_1_V(reg_q_i[5][1][1]),
.q_i_5_1_2_V(reg_q_i[5][1][2]),
.q_i_5_2_0_V(reg_q_i[5][2][0]),
.q_i_5_2_1_V(reg_q_i[5][2][1]),
.q_i_5_2_2_V(reg_q_i[5][2][2]),
.q_i_5_3_0_V(reg_q_i[5][3][0]),
.q_i_5_3_1_V(reg_q_i[5][3][1]),
.q_i_5_3_2_V(reg_q_i[5][3][2]),
.q_i_5_4_0_V(reg_q_i[5][4][0]),
.q_i_5_4_1_V(reg_q_i[5][4][1]),
.q_i_5_4_2_V(reg_q_i[5][4][2]),
.q_i_5_5_0_V(reg_q_i[5][5][0]),
.q_i_5_5_1_V(reg_q_i[5][5][1]),
.q_i_5_5_2_V(reg_q_i[5][5][2]),
.q_i_5_6_0_V(reg_q_i[5][6][0]),
.q_i_5_6_1_V(reg_q_i[5][6][1]),
.q_i_5_6_2_V(reg_q_i[5][6][2]),
.q_i_5_7_0_V(reg_q_i[5][7][0]),
.q_i_5_7_1_V(reg_q_i[5][7][1]),
.q_i_5_7_2_V(reg_q_i[5][7][2]),
.q_i_5_8_0_V(reg_q_i[5][8][0]),
.q_i_5_8_1_V(reg_q_i[5][8][1]),
.q_i_5_8_2_V(reg_q_i[5][8][2]),
.q_i_6_0_0_V(reg_q_i[6][0][0]),
.q_i_6_0_1_V(reg_q_i[6][0][1]),
.q_i_6_0_2_V(reg_q_i[6][0][2]),
.q_i_6_1_0_V(reg_q_i[6][1][0]),
.q_i_6_1_1_V(reg_q_i[6][1][1]),
.q_i_6_1_2_V(reg_q_i[6][1][2]),
.q_i_6_2_0_V(reg_q_i[6][2][0]),
.q_i_6_2_1_V(reg_q_i[6][2][1]),
.q_i_6_2_2_V(reg_q_i[6][2][2]),
.q_i_6_3_0_V(reg_q_i[6][3][0]),
.q_i_6_3_1_V(reg_q_i[6][3][1]),
.q_i_6_3_2_V(reg_q_i[6][3][2]),
.q_i_6_4_0_V(reg_q_i[6][4][0]),
.q_i_6_4_1_V(reg_q_i[6][4][1]),
.q_i_6_4_2_V(reg_q_i[6][4][2]),
.q_i_6_5_0_V(reg_q_i[6][5][0]),
.q_i_6_5_1_V(reg_q_i[6][5][1]),
.q_i_6_5_2_V(reg_q_i[6][5][2]),
.q_i_6_6_0_V(reg_q_i[6][6][0]),
.q_i_6_6_1_V(reg_q_i[6][6][1]),
.q_i_6_6_2_V(reg_q_i[6][6][2]),
.q_i_6_7_0_V(reg_q_i[6][7][0]),
.q_i_6_7_1_V(reg_q_i[6][7][1]),
.q_i_6_7_2_V(reg_q_i[6][7][2]),
.q_i_6_8_0_V(reg_q_i[6][8][0]),
.q_i_6_8_1_V(reg_q_i[6][8][1]),
.q_i_6_8_2_V(reg_q_i[6][8][2]),
.q_i_7_0_0_V(reg_q_i[7][0][0]),
.q_i_7_0_1_V(reg_q_i[7][0][1]),
.q_i_7_0_2_V(reg_q_i[7][0][2]),
.q_i_7_1_0_V(reg_q_i[7][1][0]),
.q_i_7_1_1_V(reg_q_i[7][1][1]),
.q_i_7_1_2_V(reg_q_i[7][1][2]),
.q_i_7_2_0_V(reg_q_i[7][2][0]),
.q_i_7_2_1_V(reg_q_i[7][2][1]),
.q_i_7_2_2_V(reg_q_i[7][2][2]),
.q_i_7_3_0_V(reg_q_i[7][3][0]),
.q_i_7_3_1_V(reg_q_i[7][3][1]),
.q_i_7_3_2_V(reg_q_i[7][3][2]),
.q_i_7_4_0_V(reg_q_i[7][4][0]),
.q_i_7_4_1_V(reg_q_i[7][4][1]),
.q_i_7_4_2_V(reg_q_i[7][4][2]),
.q_i_7_5_0_V(reg_q_i[7][5][0]),
.q_i_7_5_1_V(reg_q_i[7][5][1]),
.q_i_7_5_2_V(reg_q_i[7][5][2]),
.q_i_7_6_0_V(reg_q_i[7][6][0]),
.q_i_7_6_1_V(reg_q_i[7][6][1]),
.q_i_7_6_2_V(reg_q_i[7][6][2]),
.q_i_7_7_0_V(reg_q_i[7][7][0]),
.q_i_7_7_1_V(reg_q_i[7][7][1]),
.q_i_7_7_2_V(reg_q_i[7][7][2]),
.q_i_7_8_0_V(reg_q_i[7][8][0]),
.q_i_7_8_1_V(reg_q_i[7][8][1]),
.q_i_7_8_2_V(reg_q_i[7][8][2]),
.q_i_8_0_0_V(reg_q_i[8][0][0]),
.q_i_8_0_1_V(reg_q_i[8][0][1]),
.q_i_8_0_2_V(reg_q_i[8][0][2]),
.q_i_8_1_0_V(reg_q_i[8][1][0]),
.q_i_8_1_1_V(reg_q_i[8][1][1]),
.q_i_8_1_2_V(reg_q_i[8][1][2]),
.q_i_8_2_0_V(reg_q_i[8][2][0]),
.q_i_8_2_1_V(reg_q_i[8][2][1]),
.q_i_8_2_2_V(reg_q_i[8][2][2]),
.q_i_8_3_0_V(reg_q_i[8][3][0]),
.q_i_8_3_1_V(reg_q_i[8][3][1]),
.q_i_8_3_2_V(reg_q_i[8][3][2]),
.q_i_8_4_0_V(reg_q_i[8][4][0]),
.q_i_8_4_1_V(reg_q_i[8][4][1]),
.q_i_8_4_2_V(reg_q_i[8][4][2]),
.q_i_8_5_0_V(reg_q_i[8][5][0]),
.q_i_8_5_1_V(reg_q_i[8][5][1]),
.q_i_8_5_2_V(reg_q_i[8][5][2]),
.q_i_8_6_0_V(reg_q_i[8][6][0]),
.q_i_8_6_1_V(reg_q_i[8][6][1]),
.q_i_8_6_2_V(reg_q_i[8][6][2]),
.q_i_8_7_0_V(reg_q_i[8][7][0]),
.q_i_8_7_1_V(reg_q_i[8][7][1]),
.q_i_8_7_2_V(reg_q_i[8][7][2]),
.q_i_8_8_0_V(reg_q_i[8][8][0]),
.q_i_8_8_1_V(reg_q_i[8][8][1]),
.q_i_8_8_2_V(reg_q_i[8][8][2]),
.q_i_9_0_0_V(reg_q_i[9][0][0]),
.q_i_9_0_1_V(reg_q_i[9][0][1]),
.q_i_9_0_2_V(reg_q_i[9][0][2]),
.q_i_9_1_0_V(reg_q_i[9][1][0]),
.q_i_9_1_1_V(reg_q_i[9][1][1]),
.q_i_9_1_2_V(reg_q_i[9][1][2]),
.q_i_9_2_0_V(reg_q_i[9][2][0]),
.q_i_9_2_1_V(reg_q_i[9][2][1]),
.q_i_9_2_2_V(reg_q_i[9][2][2]),
.q_i_9_3_0_V(reg_q_i[9][3][0]),
.q_i_9_3_1_V(reg_q_i[9][3][1]),
.q_i_9_3_2_V(reg_q_i[9][3][2]),
.q_i_9_4_0_V(reg_q_i[9][4][0]),
.q_i_9_4_1_V(reg_q_i[9][4][1]),
.q_i_9_4_2_V(reg_q_i[9][4][2]),
.q_i_9_5_0_V(reg_q_i[9][5][0]),
.q_i_9_5_1_V(reg_q_i[9][5][1]),
.q_i_9_5_2_V(reg_q_i[9][5][2]),
.q_i_9_6_0_V(reg_q_i[9][6][0]),
.q_i_9_6_1_V(reg_q_i[9][6][1]),
.q_i_9_6_2_V(reg_q_i[9][6][2]),
.q_i_9_7_0_V(reg_q_i[9][7][0]),
.q_i_9_7_1_V(reg_q_i[9][7][1]),
.q_i_9_7_2_V(reg_q_i[9][7][2]),
.q_i_9_8_0_V(reg_q_i[9][8][0]),
.q_i_9_8_1_V(reg_q_i[9][8][1]),
.q_i_9_8_2_V(reg_q_i[9][8][2]),
.q_i_10_0_0_V(reg_q_i[10][0][0]),
.q_i_10_0_1_V(reg_q_i[10][0][1]),
.q_i_10_0_2_V(reg_q_i[10][0][2]),
.q_i_10_1_0_V(reg_q_i[10][1][0]),
.q_i_10_1_1_V(reg_q_i[10][1][1]),
.q_i_10_1_2_V(reg_q_i[10][1][2]),
.q_i_10_2_0_V(reg_q_i[10][2][0]),
.q_i_10_2_1_V(reg_q_i[10][2][1]),
.q_i_10_2_2_V(reg_q_i[10][2][2]),
.q_i_10_3_0_V(reg_q_i[10][3][0]),
.q_i_10_3_1_V(reg_q_i[10][3][1]),
.q_i_10_3_2_V(reg_q_i[10][3][2]),
.q_i_10_4_0_V(reg_q_i[10][4][0]),
.q_i_10_4_1_V(reg_q_i[10][4][1]),
.q_i_10_4_2_V(reg_q_i[10][4][2]),
.q_i_10_5_0_V(reg_q_i[10][5][0]),
.q_i_10_5_1_V(reg_q_i[10][5][1]),
.q_i_10_5_2_V(reg_q_i[10][5][2]),
.q_i_10_6_0_V(reg_q_i[10][6][0]),
.q_i_10_6_1_V(reg_q_i[10][6][1]),
.q_i_10_6_2_V(reg_q_i[10][6][2]),
.q_i_10_7_0_V(reg_q_i[10][7][0]),
.q_i_10_7_1_V(reg_q_i[10][7][1]),
.q_i_10_7_2_V(reg_q_i[10][7][2]),
.q_i_10_8_0_V(reg_q_i[10][8][0]),
.q_i_10_8_1_V(reg_q_i[10][8][1]),
.q_i_10_8_2_V(reg_q_i[10][8][2]),
.q_i_11_0_0_V(reg_q_i[11][0][0]),
.q_i_11_0_1_V(reg_q_i[11][0][1]),
.q_i_11_0_2_V(reg_q_i[11][0][2]),
.q_i_11_1_0_V(reg_q_i[11][1][0]),
.q_i_11_1_1_V(reg_q_i[11][1][1]),
.q_i_11_1_2_V(reg_q_i[11][1][2]),
.q_i_11_2_0_V(reg_q_i[11][2][0]),
.q_i_11_2_1_V(reg_q_i[11][2][1]),
.q_i_11_2_2_V(reg_q_i[11][2][2]),
.q_i_11_3_0_V(reg_q_i[11][3][0]),
.q_i_11_3_1_V(reg_q_i[11][3][1]),
.q_i_11_3_2_V(reg_q_i[11][3][2]),
.q_i_11_4_0_V(reg_q_i[11][4][0]),
.q_i_11_4_1_V(reg_q_i[11][4][1]),
.q_i_11_4_2_V(reg_q_i[11][4][2]),
.q_i_11_5_0_V(reg_q_i[11][5][0]),
.q_i_11_5_1_V(reg_q_i[11][5][1]),
.q_i_11_5_2_V(reg_q_i[11][5][2]),
.q_i_11_6_0_V(reg_q_i[11][6][0]),
.q_i_11_6_1_V(reg_q_i[11][6][1]),
.q_i_11_6_2_V(reg_q_i[11][6][2]),
.q_i_11_7_0_V(reg_q_i[11][7][0]),
.q_i_11_7_1_V(reg_q_i[11][7][1]),
.q_i_11_7_2_V(reg_q_i[11][7][2]),
.q_i_11_8_0_V(reg_q_i[11][8][0]),
.q_i_11_8_1_V(reg_q_i[11][8][1]),
.q_i_11_8_2_V(reg_q_i[11][8][2]),
.q_i_12_0_0_V(reg_q_i[12][0][0]),
.q_i_12_0_1_V(reg_q_i[12][0][1]),
.q_i_12_0_2_V(reg_q_i[12][0][2]),
.q_i_12_1_0_V(reg_q_i[12][1][0]),
.q_i_12_1_1_V(reg_q_i[12][1][1]),
.q_i_12_1_2_V(reg_q_i[12][1][2]),
.q_i_12_2_0_V(reg_q_i[12][2][0]),
.q_i_12_2_1_V(reg_q_i[12][2][1]),
.q_i_12_2_2_V(reg_q_i[12][2][2]),
.q_i_12_3_0_V(reg_q_i[12][3][0]),
.q_i_12_3_1_V(reg_q_i[12][3][1]),
.q_i_12_3_2_V(reg_q_i[12][3][2]),
.q_i_12_4_0_V(reg_q_i[12][4][0]),
.q_i_12_4_1_V(reg_q_i[12][4][1]),
.q_i_12_4_2_V(reg_q_i[12][4][2]),
.q_i_12_5_0_V(reg_q_i[12][5][0]),
.q_i_12_5_1_V(reg_q_i[12][5][1]),
.q_i_12_5_2_V(reg_q_i[12][5][2]),
.q_i_12_6_0_V(reg_q_i[12][6][0]),
.q_i_12_6_1_V(reg_q_i[12][6][1]),
.q_i_12_6_2_V(reg_q_i[12][6][2]),
.q_i_12_7_0_V(reg_q_i[12][7][0]),
.q_i_12_7_1_V(reg_q_i[12][7][1]),
.q_i_12_7_2_V(reg_q_i[12][7][2]),
.q_i_12_8_0_V(reg_q_i[12][8][0]),
.q_i_12_8_1_V(reg_q_i[12][8][1]),
.q_i_12_8_2_V(reg_q_i[12][8][2]),
.cpatr_i_0_0_0_V(reg_cpatr_i[0][0][0]),
.cpatr_i_0_0_1_V(reg_cpatr_i[0][0][1]),
.cpatr_i_0_1_0_V(reg_cpatr_i[0][1][0]),
.cpatr_i_0_1_1_V(reg_cpatr_i[0][1][1]),
.cpatr_i_0_2_0_V(reg_cpatr_i[0][2][0]),
.cpatr_i_0_2_1_V(reg_cpatr_i[0][2][1]),
.cpatr_i_0_3_0_V(reg_cpatr_i[0][3][0]),
.cpatr_i_0_3_1_V(reg_cpatr_i[0][3][1]),
.cpatr_i_0_4_0_V(reg_cpatr_i[0][4][0]),
.cpatr_i_0_4_1_V(reg_cpatr_i[0][4][1]),
.cpatr_i_0_5_0_V(reg_cpatr_i[0][5][0]),
.cpatr_i_0_5_1_V(reg_cpatr_i[0][5][1]),
.cpatr_i_0_6_0_V(reg_cpatr_i[0][6][0]),
.cpatr_i_0_6_1_V(reg_cpatr_i[0][6][1]),
.cpatr_i_0_7_0_V(reg_cpatr_i[0][7][0]),
.cpatr_i_0_7_1_V(reg_cpatr_i[0][7][1]),
.cpatr_i_0_8_0_V(reg_cpatr_i[0][8][0]),
.cpatr_i_0_8_1_V(reg_cpatr_i[0][8][1]),
.cpatr_i_1_0_0_V(reg_cpatr_i[1][0][0]),
.cpatr_i_1_0_1_V(reg_cpatr_i[1][0][1]),
.cpatr_i_1_1_0_V(reg_cpatr_i[1][1][0]),
.cpatr_i_1_1_1_V(reg_cpatr_i[1][1][1]),
.cpatr_i_1_2_0_V(reg_cpatr_i[1][2][0]),
.cpatr_i_1_2_1_V(reg_cpatr_i[1][2][1]),
.cpatr_i_1_3_0_V(reg_cpatr_i[1][3][0]),
.cpatr_i_1_3_1_V(reg_cpatr_i[1][3][1]),
.cpatr_i_1_4_0_V(reg_cpatr_i[1][4][0]),
.cpatr_i_1_4_1_V(reg_cpatr_i[1][4][1]),
.cpatr_i_1_5_0_V(reg_cpatr_i[1][5][0]),
.cpatr_i_1_5_1_V(reg_cpatr_i[1][5][1]),
.cpatr_i_1_6_0_V(reg_cpatr_i[1][6][0]),
.cpatr_i_1_6_1_V(reg_cpatr_i[1][6][1]),
.cpatr_i_1_7_0_V(reg_cpatr_i[1][7][0]),
.cpatr_i_1_7_1_V(reg_cpatr_i[1][7][1]),
.cpatr_i_1_8_0_V(reg_cpatr_i[1][8][0]),
.cpatr_i_1_8_1_V(reg_cpatr_i[1][8][1]),
.cpatr_i_2_0_0_V(reg_cpatr_i[2][0][0]),
.cpatr_i_2_0_1_V(reg_cpatr_i[2][0][1]),
.cpatr_i_2_1_0_V(reg_cpatr_i[2][1][0]),
.cpatr_i_2_1_1_V(reg_cpatr_i[2][1][1]),
.cpatr_i_2_2_0_V(reg_cpatr_i[2][2][0]),
.cpatr_i_2_2_1_V(reg_cpatr_i[2][2][1]),
.cpatr_i_2_3_0_V(reg_cpatr_i[2][3][0]),
.cpatr_i_2_3_1_V(reg_cpatr_i[2][3][1]),
.cpatr_i_2_4_0_V(reg_cpatr_i[2][4][0]),
.cpatr_i_2_4_1_V(reg_cpatr_i[2][4][1]),
.cpatr_i_2_5_0_V(reg_cpatr_i[2][5][0]),
.cpatr_i_2_5_1_V(reg_cpatr_i[2][5][1]),
.cpatr_i_2_6_0_V(reg_cpatr_i[2][6][0]),
.cpatr_i_2_6_1_V(reg_cpatr_i[2][6][1]),
.cpatr_i_2_7_0_V(reg_cpatr_i[2][7][0]),
.cpatr_i_2_7_1_V(reg_cpatr_i[2][7][1]),
.cpatr_i_2_8_0_V(reg_cpatr_i[2][8][0]),
.cpatr_i_2_8_1_V(reg_cpatr_i[2][8][1]),
.cpatr_i_3_0_0_V(reg_cpatr_i[3][0][0]),
.cpatr_i_3_0_1_V(reg_cpatr_i[3][0][1]),
.cpatr_i_3_1_0_V(reg_cpatr_i[3][1][0]),
.cpatr_i_3_1_1_V(reg_cpatr_i[3][1][1]),
.cpatr_i_3_2_0_V(reg_cpatr_i[3][2][0]),
.cpatr_i_3_2_1_V(reg_cpatr_i[3][2][1]),
.cpatr_i_3_3_0_V(reg_cpatr_i[3][3][0]),
.cpatr_i_3_3_1_V(reg_cpatr_i[3][3][1]),
.cpatr_i_3_4_0_V(reg_cpatr_i[3][4][0]),
.cpatr_i_3_4_1_V(reg_cpatr_i[3][4][1]),
.cpatr_i_3_5_0_V(reg_cpatr_i[3][5][0]),
.cpatr_i_3_5_1_V(reg_cpatr_i[3][5][1]),
.cpatr_i_3_6_0_V(reg_cpatr_i[3][6][0]),
.cpatr_i_3_6_1_V(reg_cpatr_i[3][6][1]),
.cpatr_i_3_7_0_V(reg_cpatr_i[3][7][0]),
.cpatr_i_3_7_1_V(reg_cpatr_i[3][7][1]),
.cpatr_i_3_8_0_V(reg_cpatr_i[3][8][0]),
.cpatr_i_3_8_1_V(reg_cpatr_i[3][8][1]),
.cpatr_i_4_0_0_V(reg_cpatr_i[4][0][0]),
.cpatr_i_4_0_1_V(reg_cpatr_i[4][0][1]),
.cpatr_i_4_1_0_V(reg_cpatr_i[4][1][0]),
.cpatr_i_4_1_1_V(reg_cpatr_i[4][1][1]),
.cpatr_i_4_2_0_V(reg_cpatr_i[4][2][0]),
.cpatr_i_4_2_1_V(reg_cpatr_i[4][2][1]),
.cpatr_i_4_3_0_V(reg_cpatr_i[4][3][0]),
.cpatr_i_4_3_1_V(reg_cpatr_i[4][3][1]),
.cpatr_i_4_4_0_V(reg_cpatr_i[4][4][0]),
.cpatr_i_4_4_1_V(reg_cpatr_i[4][4][1]),
.cpatr_i_4_5_0_V(reg_cpatr_i[4][5][0]),
.cpatr_i_4_5_1_V(reg_cpatr_i[4][5][1]),
.cpatr_i_4_6_0_V(reg_cpatr_i[4][6][0]),
.cpatr_i_4_6_1_V(reg_cpatr_i[4][6][1]),
.cpatr_i_4_7_0_V(reg_cpatr_i[4][7][0]),
.cpatr_i_4_7_1_V(reg_cpatr_i[4][7][1]),
.cpatr_i_4_8_0_V(reg_cpatr_i[4][8][0]),
.cpatr_i_4_8_1_V(reg_cpatr_i[4][8][1]),
.cpatr_i_5_0_0_V(reg_cpatr_i[5][0][0]),
.cpatr_i_5_0_1_V(reg_cpatr_i[5][0][1]),
.cpatr_i_5_1_0_V(reg_cpatr_i[5][1][0]),
.cpatr_i_5_1_1_V(reg_cpatr_i[5][1][1]),
.cpatr_i_5_2_0_V(reg_cpatr_i[5][2][0]),
.cpatr_i_5_2_1_V(reg_cpatr_i[5][2][1]),
.cpatr_i_5_3_0_V(reg_cpatr_i[5][3][0]),
.cpatr_i_5_3_1_V(reg_cpatr_i[5][3][1]),
.cpatr_i_5_4_0_V(reg_cpatr_i[5][4][0]),
.cpatr_i_5_4_1_V(reg_cpatr_i[5][4][1]),
.cpatr_i_5_5_0_V(reg_cpatr_i[5][5][0]),
.cpatr_i_5_5_1_V(reg_cpatr_i[5][5][1]),
.cpatr_i_5_6_0_V(reg_cpatr_i[5][6][0]),
.cpatr_i_5_6_1_V(reg_cpatr_i[5][6][1]),
.cpatr_i_5_7_0_V(reg_cpatr_i[5][7][0]),
.cpatr_i_5_7_1_V(reg_cpatr_i[5][7][1]),
.cpatr_i_5_8_0_V(reg_cpatr_i[5][8][0]),
.cpatr_i_5_8_1_V(reg_cpatr_i[5][8][1]),
.ph_i_0_0_0_V(reg_ph_i[0][0][0]),
.ph_i_0_0_1_V(reg_ph_i[0][0][1]),
.ph_i_0_1_0_V(reg_ph_i[0][1][0]),
.ph_i_0_1_1_V(reg_ph_i[0][1][1]),
.ph_i_0_2_0_V(reg_ph_i[0][2][0]),
.ph_i_0_2_1_V(reg_ph_i[0][2][1]),
.ph_i_0_3_0_V(reg_ph_i[0][3][0]),
.ph_i_0_3_1_V(reg_ph_i[0][3][1]),
.ph_i_0_4_0_V(reg_ph_i[0][4][0]),
.ph_i_0_4_1_V(reg_ph_i[0][4][1]),
.ph_i_0_5_0_V(reg_ph_i[0][5][0]),
.ph_i_0_5_1_V(reg_ph_i[0][5][1]),
.ph_i_0_6_0_V(reg_ph_i[0][6][0]),
.ph_i_0_6_1_V(reg_ph_i[0][6][1]),
.ph_i_0_7_0_V(reg_ph_i[0][7][0]),
.ph_i_0_7_1_V(reg_ph_i[0][7][1]),
.ph_i_0_8_0_V(reg_ph_i[0][8][0]),
.ph_i_0_8_1_V(reg_ph_i[0][8][1]),
.ph_i_1_0_0_V(reg_ph_i[1][0][0]),
.ph_i_1_0_1_V(reg_ph_i[1][0][1]),
.ph_i_1_1_0_V(reg_ph_i[1][1][0]),
.ph_i_1_1_1_V(reg_ph_i[1][1][1]),
.ph_i_1_2_0_V(reg_ph_i[1][2][0]),
.ph_i_1_2_1_V(reg_ph_i[1][2][1]),
.ph_i_1_3_0_V(reg_ph_i[1][3][0]),
.ph_i_1_3_1_V(reg_ph_i[1][3][1]),
.ph_i_1_4_0_V(reg_ph_i[1][4][0]),
.ph_i_1_4_1_V(reg_ph_i[1][4][1]),
.ph_i_1_5_0_V(reg_ph_i[1][5][0]),
.ph_i_1_5_1_V(reg_ph_i[1][5][1]),
.ph_i_1_6_0_V(reg_ph_i[1][6][0]),
.ph_i_1_6_1_V(reg_ph_i[1][6][1]),
.ph_i_1_7_0_V(reg_ph_i[1][7][0]),
.ph_i_1_7_1_V(reg_ph_i[1][7][1]),
.ph_i_1_8_0_V(reg_ph_i[1][8][0]),
.ph_i_1_8_1_V(reg_ph_i[1][8][1]),
.ph_i_2_0_0_V(reg_ph_i[2][0][0]),
.ph_i_2_0_1_V(reg_ph_i[2][0][1]),
.ph_i_2_1_0_V(reg_ph_i[2][1][0]),
.ph_i_2_1_1_V(reg_ph_i[2][1][1]),
.ph_i_2_2_0_V(reg_ph_i[2][2][0]),
.ph_i_2_2_1_V(reg_ph_i[2][2][1]),
.ph_i_2_3_0_V(reg_ph_i[2][3][0]),
.ph_i_2_3_1_V(reg_ph_i[2][3][1]),
.ph_i_2_4_0_V(reg_ph_i[2][4][0]),
.ph_i_2_4_1_V(reg_ph_i[2][4][1]),
.ph_i_2_5_0_V(reg_ph_i[2][5][0]),
.ph_i_2_5_1_V(reg_ph_i[2][5][1]),
.ph_i_2_6_0_V(reg_ph_i[2][6][0]),
.ph_i_2_6_1_V(reg_ph_i[2][6][1]),
.ph_i_2_7_0_V(reg_ph_i[2][7][0]),
.ph_i_2_7_1_V(reg_ph_i[2][7][1]),
.ph_i_2_8_0_V(reg_ph_i[2][8][0]),
.ph_i_2_8_1_V(reg_ph_i[2][8][1]),
.ph_i_3_0_0_V(reg_ph_i[3][0][0]),
.ph_i_3_0_1_V(reg_ph_i[3][0][1]),
.ph_i_3_1_0_V(reg_ph_i[3][1][0]),
.ph_i_3_1_1_V(reg_ph_i[3][1][1]),
.ph_i_3_2_0_V(reg_ph_i[3][2][0]),
.ph_i_3_2_1_V(reg_ph_i[3][2][1]),
.ph_i_3_3_0_V(reg_ph_i[3][3][0]),
.ph_i_3_3_1_V(reg_ph_i[3][3][1]),
.ph_i_3_4_0_V(reg_ph_i[3][4][0]),
.ph_i_3_4_1_V(reg_ph_i[3][4][1]),
.ph_i_3_5_0_V(reg_ph_i[3][5][0]),
.ph_i_3_5_1_V(reg_ph_i[3][5][1]),
.ph_i_3_6_0_V(reg_ph_i[3][6][0]),
.ph_i_3_6_1_V(reg_ph_i[3][6][1]),
.ph_i_3_7_0_V(reg_ph_i[3][7][0]),
.ph_i_3_7_1_V(reg_ph_i[3][7][1]),
.ph_i_3_8_0_V(reg_ph_i[3][8][0]),
.ph_i_3_8_1_V(reg_ph_i[3][8][1]),
.ph_i_4_0_0_V(reg_ph_i[4][0][0]),
.ph_i_4_0_1_V(reg_ph_i[4][0][1]),
.ph_i_4_1_0_V(reg_ph_i[4][1][0]),
.ph_i_4_1_1_V(reg_ph_i[4][1][1]),
.ph_i_4_2_0_V(reg_ph_i[4][2][0]),
.ph_i_4_2_1_V(reg_ph_i[4][2][1]),
.ph_i_4_3_0_V(reg_ph_i[4][3][0]),
.ph_i_4_3_1_V(reg_ph_i[4][3][1]),
.ph_i_4_4_0_V(reg_ph_i[4][4][0]),
.ph_i_4_4_1_V(reg_ph_i[4][4][1]),
.ph_i_4_5_0_V(reg_ph_i[4][5][0]),
.ph_i_4_5_1_V(reg_ph_i[4][5][1]),
.ph_i_4_6_0_V(reg_ph_i[4][6][0]),
.ph_i_4_6_1_V(reg_ph_i[4][6][1]),
.ph_i_4_7_0_V(reg_ph_i[4][7][0]),
.ph_i_4_7_1_V(reg_ph_i[4][7][1]),
.ph_i_4_8_0_V(reg_ph_i[4][8][0]),
.ph_i_4_8_1_V(reg_ph_i[4][8][1]),
.ph_i_5_0_0_V(reg_ph_i[5][0][0]),
.ph_i_5_0_1_V(reg_ph_i[5][0][1]),
.ph_i_5_1_0_V(reg_ph_i[5][1][0]),
.ph_i_5_1_1_V(reg_ph_i[5][1][1]),
.ph_i_5_2_0_V(reg_ph_i[5][2][0]),
.ph_i_5_2_1_V(reg_ph_i[5][2][1]),
.ph_i_5_3_0_V(reg_ph_i[5][3][0]),
.ph_i_5_3_1_V(reg_ph_i[5][3][1]),
.ph_i_5_4_0_V(reg_ph_i[5][4][0]),
.ph_i_5_4_1_V(reg_ph_i[5][4][1]),
.ph_i_5_5_0_V(reg_ph_i[5][5][0]),
.ph_i_5_5_1_V(reg_ph_i[5][5][1]),
.ph_i_5_6_0_V(reg_ph_i[5][6][0]),
.ph_i_5_6_1_V(reg_ph_i[5][6][1]),
.ph_i_5_7_0_V(reg_ph_i[5][7][0]),
.ph_i_5_7_1_V(reg_ph_i[5][7][1]),
.ph_i_5_8_0_V(reg_ph_i[5][8][0]),
.ph_i_5_8_1_V(reg_ph_i[5][8][1]),
.th11_i_0_0_0_V(reg_th11_i[0][0][0]),
.th11_i_0_0_1_V(reg_th11_i[0][0][1]),
.th11_i_0_1_0_V(reg_th11_i[0][1][0]),
.th11_i_0_1_1_V(reg_th11_i[0][1][1]),
.th11_i_0_2_0_V(reg_th11_i[0][2][0]),
.th11_i_0_2_1_V(reg_th11_i[0][2][1]),
.th11_i_0_3_0_V(reg_th11_i[0][3][0]),
.th11_i_0_3_1_V(reg_th11_i[0][3][1]),
.th11_i_0_4_0_V(reg_th11_i[0][4][0]),
.th11_i_0_4_1_V(reg_th11_i[0][4][1]),
.th11_i_0_5_0_V(reg_th11_i[0][5][0]),
.th11_i_0_5_1_V(reg_th11_i[0][5][1]),
.th11_i_0_6_0_V(reg_th11_i[0][6][0]),
.th11_i_0_6_1_V(reg_th11_i[0][6][1]),
.th11_i_0_7_0_V(reg_th11_i[0][7][0]),
.th11_i_0_7_1_V(reg_th11_i[0][7][1]),
.th11_i_0_8_0_V(reg_th11_i[0][8][0]),
.th11_i_0_8_1_V(reg_th11_i[0][8][1]),
.th11_i_1_0_0_V(reg_th11_i[1][0][0]),
.th11_i_1_0_1_V(reg_th11_i[1][0][1]),
.th11_i_1_1_0_V(reg_th11_i[1][1][0]),
.th11_i_1_1_1_V(reg_th11_i[1][1][1]),
.th11_i_1_2_0_V(reg_th11_i[1][2][0]),
.th11_i_1_2_1_V(reg_th11_i[1][2][1]),
.th11_i_1_3_0_V(reg_th11_i[1][3][0]),
.th11_i_1_3_1_V(reg_th11_i[1][3][1]),
.th11_i_1_4_0_V(reg_th11_i[1][4][0]),
.th11_i_1_4_1_V(reg_th11_i[1][4][1]),
.th11_i_1_5_0_V(reg_th11_i[1][5][0]),
.th11_i_1_5_1_V(reg_th11_i[1][5][1]),
.th11_i_1_6_0_V(reg_th11_i[1][6][0]),
.th11_i_1_6_1_V(reg_th11_i[1][6][1]),
.th11_i_1_7_0_V(reg_th11_i[1][7][0]),
.th11_i_1_7_1_V(reg_th11_i[1][7][1]),
.th11_i_1_8_0_V(reg_th11_i[1][8][0]),
.th11_i_1_8_1_V(reg_th11_i[1][8][1]),
.th11_i_2_0_0_V(reg_th11_i[2][0][0]),
.th11_i_2_0_1_V(reg_th11_i[2][0][1]),
.th11_i_2_1_0_V(reg_th11_i[2][1][0]),
.th11_i_2_1_1_V(reg_th11_i[2][1][1]),
.th11_i_2_2_0_V(reg_th11_i[2][2][0]),
.th11_i_2_2_1_V(reg_th11_i[2][2][1]),
.th11_i_2_3_0_V(reg_th11_i[2][3][0]),
.th11_i_2_3_1_V(reg_th11_i[2][3][1]),
.th11_i_2_4_0_V(reg_th11_i[2][4][0]),
.th11_i_2_4_1_V(reg_th11_i[2][4][1]),
.th11_i_2_5_0_V(reg_th11_i[2][5][0]),
.th11_i_2_5_1_V(reg_th11_i[2][5][1]),
.th11_i_2_6_0_V(reg_th11_i[2][6][0]),
.th11_i_2_6_1_V(reg_th11_i[2][6][1]),
.th11_i_2_7_0_V(reg_th11_i[2][7][0]),
.th11_i_2_7_1_V(reg_th11_i[2][7][1]),
.th11_i_2_8_0_V(reg_th11_i[2][8][0]),
.th11_i_2_8_1_V(reg_th11_i[2][8][1]),
.th11_i_3_0_0_V(reg_th11_i[3][0][0]),
.th11_i_3_0_1_V(reg_th11_i[3][0][1]),
.th11_i_3_1_0_V(reg_th11_i[3][1][0]),
.th11_i_3_1_1_V(reg_th11_i[3][1][1]),
.th11_i_3_2_0_V(reg_th11_i[3][2][0]),
.th11_i_3_2_1_V(reg_th11_i[3][2][1]),
.th11_i_3_3_0_V(reg_th11_i[3][3][0]),
.th11_i_3_3_1_V(reg_th11_i[3][3][1]),
.th11_i_3_4_0_V(reg_th11_i[3][4][0]),
.th11_i_3_4_1_V(reg_th11_i[3][4][1]),
.th11_i_3_5_0_V(reg_th11_i[3][5][0]),
.th11_i_3_5_1_V(reg_th11_i[3][5][1]),
.th11_i_3_6_0_V(reg_th11_i[3][6][0]),
.th11_i_3_6_1_V(reg_th11_i[3][6][1]),
.th11_i_3_7_0_V(reg_th11_i[3][7][0]),
.th11_i_3_7_1_V(reg_th11_i[3][7][1]),
.th11_i_3_8_0_V(reg_th11_i[3][8][0]),
.th11_i_3_8_1_V(reg_th11_i[3][8][1]),
.th11_i_4_0_0_V(reg_th11_i[4][0][0]),
.th11_i_4_0_1_V(reg_th11_i[4][0][1]),
.th11_i_4_1_0_V(reg_th11_i[4][1][0]),
.th11_i_4_1_1_V(reg_th11_i[4][1][1]),
.th11_i_4_2_0_V(reg_th11_i[4][2][0]),
.th11_i_4_2_1_V(reg_th11_i[4][2][1]),
.th11_i_4_3_0_V(reg_th11_i[4][3][0]),
.th11_i_4_3_1_V(reg_th11_i[4][3][1]),
.th11_i_4_4_0_V(reg_th11_i[4][4][0]),
.th11_i_4_4_1_V(reg_th11_i[4][4][1]),
.th11_i_4_5_0_V(reg_th11_i[4][5][0]),
.th11_i_4_5_1_V(reg_th11_i[4][5][1]),
.th11_i_4_6_0_V(reg_th11_i[4][6][0]),
.th11_i_4_6_1_V(reg_th11_i[4][6][1]),
.th11_i_4_7_0_V(reg_th11_i[4][7][0]),
.th11_i_4_7_1_V(reg_th11_i[4][7][1]),
.th11_i_4_8_0_V(reg_th11_i[4][8][0]),
.th11_i_4_8_1_V(reg_th11_i[4][8][1]),
.th11_i_5_0_0_V(reg_th11_i[5][0][0]),
.th11_i_5_0_1_V(reg_th11_i[5][0][1]),
.th11_i_5_1_0_V(reg_th11_i[5][1][0]),
.th11_i_5_1_1_V(reg_th11_i[5][1][1]),
.th11_i_5_2_0_V(reg_th11_i[5][2][0]),
.th11_i_5_2_1_V(reg_th11_i[5][2][1]),
.th11_i_5_3_0_V(reg_th11_i[5][3][0]),
.th11_i_5_3_1_V(reg_th11_i[5][3][1]),
.th11_i_5_4_0_V(reg_th11_i[5][4][0]),
.th11_i_5_4_1_V(reg_th11_i[5][4][1]),
.th11_i_5_5_0_V(reg_th11_i[5][5][0]),
.th11_i_5_5_1_V(reg_th11_i[5][5][1]),
.th11_i_5_6_0_V(reg_th11_i[5][6][0]),
.th11_i_5_6_1_V(reg_th11_i[5][6][1]),
.th11_i_5_7_0_V(reg_th11_i[5][7][0]),
.th11_i_5_7_1_V(reg_th11_i[5][7][1]),
.th11_i_5_8_0_V(reg_th11_i[5][8][0]),
.th11_i_5_8_1_V(reg_th11_i[5][8][1]),
.th_i_0_0_0_V(reg_th_i[0][0][0]),
.th_i_0_0_1_V(reg_th_i[0][0][1]),
.th_i_0_0_2_V(reg_th_i[0][0][2]),
.th_i_0_0_3_V(reg_th_i[0][0][3]),
.th_i_0_1_0_V(reg_th_i[0][1][0]),
.th_i_0_1_1_V(reg_th_i[0][1][1]),
.th_i_0_1_2_V(reg_th_i[0][1][2]),
.th_i_0_1_3_V(reg_th_i[0][1][3]),
.th_i_0_2_0_V(reg_th_i[0][2][0]),
.th_i_0_2_1_V(reg_th_i[0][2][1]),
.th_i_0_2_2_V(reg_th_i[0][2][2]),
.th_i_0_2_3_V(reg_th_i[0][2][3]),
.th_i_1_0_0_V(reg_th_i[1][0][0]),
.th_i_1_0_1_V(reg_th_i[1][0][1]),
.th_i_1_0_2_V(reg_th_i[1][0][2]),
.th_i_1_0_3_V(reg_th_i[1][0][3]),
.th_i_1_1_0_V(reg_th_i[1][1][0]),
.th_i_1_1_1_V(reg_th_i[1][1][1]),
.th_i_1_1_2_V(reg_th_i[1][1][2]),
.th_i_1_1_3_V(reg_th_i[1][1][3]),
.th_i_1_2_0_V(reg_th_i[1][2][0]),
.th_i_1_2_1_V(reg_th_i[1][2][1]),
.th_i_1_2_2_V(reg_th_i[1][2][2]),
.th_i_1_2_3_V(reg_th_i[1][2][3]),
.th_i_2_0_0_V(reg_th_i[2][0][0]),
.th_i_2_0_1_V(reg_th_i[2][0][1]),
.th_i_2_0_2_V(reg_th_i[2][0][2]),
.th_i_2_0_3_V(reg_th_i[2][0][3]),
.th_i_2_1_0_V(reg_th_i[2][1][0]),
.th_i_2_1_1_V(reg_th_i[2][1][1]),
.th_i_2_1_2_V(reg_th_i[2][1][2]),
.th_i_2_1_3_V(reg_th_i[2][1][3]),
.th_i_2_2_0_V(reg_th_i[2][2][0]),
.th_i_2_2_1_V(reg_th_i[2][2][1]),
.th_i_2_2_2_V(reg_th_i[2][2][2]),
.th_i_2_2_3_V(reg_th_i[2][2][3]),
.phzvl_i_0_0_V(reg_phzvl_i[0][0]),
.phzvl_i_0_1_V(reg_phzvl_i[0][1]),
.phzvl_i_0_2_V(reg_phzvl_i[0][2]),
.phzvl_i_0_3_V(reg_phzvl_i[0][3]),
.phzvl_i_0_4_V(reg_phzvl_i[0][4]),
.phzvl_i_0_5_V(reg_phzvl_i[0][5]),
.phzvl_i_0_6_V(reg_phzvl_i[0][6]),
.phzvl_i_0_7_V(reg_phzvl_i[0][7]),
.phzvl_i_0_8_V(reg_phzvl_i[0][8]),
.phzvl_i_1_0_V(reg_phzvl_i[1][0]),
.phzvl_i_1_1_V(reg_phzvl_i[1][1]),
.phzvl_i_1_2_V(reg_phzvl_i[1][2]),
.phzvl_i_1_3_V(reg_phzvl_i[1][3]),
.phzvl_i_1_4_V(reg_phzvl_i[1][4]),
.phzvl_i_1_5_V(reg_phzvl_i[1][5]),
.phzvl_i_1_6_V(reg_phzvl_i[1][6]),
.phzvl_i_1_7_V(reg_phzvl_i[1][7]),
.phzvl_i_1_8_V(reg_phzvl_i[1][8]),
.phzvl_i_2_0_V(reg_phzvl_i[2][0]),
.phzvl_i_2_1_V(reg_phzvl_i[2][1]),
.phzvl_i_2_2_V(reg_phzvl_i[2][2]),
.phzvl_i_2_3_V(reg_phzvl_i[2][3]),
.phzvl_i_2_4_V(reg_phzvl_i[2][4]),
.phzvl_i_2_5_V(reg_phzvl_i[2][5]),
.phzvl_i_2_6_V(reg_phzvl_i[2][6]),
.phzvl_i_2_7_V(reg_phzvl_i[2][7]),
.phzvl_i_2_8_V(reg_phzvl_i[2][8]),
.phzvl_i_3_0_V(reg_phzvl_i[3][0]),
.phzvl_i_3_1_V(reg_phzvl_i[3][1]),
.phzvl_i_3_2_V(reg_phzvl_i[3][2]),
.phzvl_i_3_3_V(reg_phzvl_i[3][3]),
.phzvl_i_3_4_V(reg_phzvl_i[3][4]),
.phzvl_i_3_5_V(reg_phzvl_i[3][5]),
.phzvl_i_3_6_V(reg_phzvl_i[3][6]),
.phzvl_i_3_7_V(reg_phzvl_i[3][7]),
.phzvl_i_3_8_V(reg_phzvl_i[3][8]),
.phzvl_i_4_0_V(reg_phzvl_i[4][0]),
.phzvl_i_4_1_V(reg_phzvl_i[4][1]),
.phzvl_i_4_2_V(reg_phzvl_i[4][2]),
.phzvl_i_4_3_V(reg_phzvl_i[4][3]),
.phzvl_i_4_4_V(reg_phzvl_i[4][4]),
.phzvl_i_4_5_V(reg_phzvl_i[4][5]),
.phzvl_i_4_6_V(reg_phzvl_i[4][6]),
.phzvl_i_4_7_V(reg_phzvl_i[4][7]),
.phzvl_i_4_8_V(reg_phzvl_i[4][8]),
.phzvl_i_5_0_V(reg_phzvl_i[5][0]),
.phzvl_i_5_1_V(reg_phzvl_i[5][1]),
.phzvl_i_5_2_V(reg_phzvl_i[5][2]),
.phzvl_i_5_3_V(reg_phzvl_i[5][3]),
.phzvl_i_5_4_V(reg_phzvl_i[5][4]),
.phzvl_i_5_5_V(reg_phzvl_i[5][5]),
.phzvl_i_5_6_V(reg_phzvl_i[5][6]),
.phzvl_i_5_7_V(reg_phzvl_i[5][7]),
.phzvl_i_5_8_V(reg_phzvl_i[5][8]),
.phzvl_i_6_0_V(reg_phzvl_i[6][0]),
.phzvl_i_6_1_V(reg_phzvl_i[6][1]),
.phzvl_i_6_2_V(reg_phzvl_i[6][2]),
.phzvl_i_6_3_V(reg_phzvl_i[6][3]),
.phzvl_i_6_4_V(reg_phzvl_i[6][4]),
.phzvl_i_6_5_V(reg_phzvl_i[6][5]),
.phzvl_i_6_6_V(reg_phzvl_i[6][6]),
.phzvl_i_6_7_V(reg_phzvl_i[6][7]),
.phzvl_i_6_8_V(reg_phzvl_i[6][8]),
.phzvl_i_7_0_V(reg_phzvl_i[7][0]),
.phzvl_i_7_1_V(reg_phzvl_i[7][1]),
.phzvl_i_7_2_V(reg_phzvl_i[7][2]),
.phzvl_i_7_3_V(reg_phzvl_i[7][3]),
.phzvl_i_7_4_V(reg_phzvl_i[7][4]),
.phzvl_i_7_5_V(reg_phzvl_i[7][5]),
.phzvl_i_7_6_V(reg_phzvl_i[7][6]),
.phzvl_i_7_7_V(reg_phzvl_i[7][7]),
.phzvl_i_7_8_V(reg_phzvl_i[7][8]),
.phzvl_i_8_0_V(reg_phzvl_i[8][0]),
.phzvl_i_8_1_V(reg_phzvl_i[8][1]),
.phzvl_i_8_2_V(reg_phzvl_i[8][2]),
.phzvl_i_8_3_V(reg_phzvl_i[8][3]),
.phzvl_i_8_4_V(reg_phzvl_i[8][4]),
.phzvl_i_8_5_V(reg_phzvl_i[8][5]),
.phzvl_i_8_6_V(reg_phzvl_i[8][6]),
.phzvl_i_8_7_V(reg_phzvl_i[8][7]),
.phzvl_i_8_8_V(reg_phzvl_i[8][8]),
.phzvl_i_9_0_V(reg_phzvl_i[9][0]),
.phzvl_i_9_1_V(reg_phzvl_i[9][1]),
.phzvl_i_9_2_V(reg_phzvl_i[9][2]),
.phzvl_i_9_3_V(reg_phzvl_i[9][3]),
.phzvl_i_9_4_V(reg_phzvl_i[9][4]),
.phzvl_i_9_5_V(reg_phzvl_i[9][5]),
.phzvl_i_9_6_V(reg_phzvl_i[9][6]),
.phzvl_i_9_7_V(reg_phzvl_i[9][7]),
.phzvl_i_9_8_V(reg_phzvl_i[9][8]),
.phzvl_i_10_0_V(reg_phzvl_i[10][0]),
.phzvl_i_10_1_V(reg_phzvl_i[10][1]),
.phzvl_i_10_2_V(reg_phzvl_i[10][2]),
.phzvl_i_10_3_V(reg_phzvl_i[10][3]),
.phzvl_i_10_4_V(reg_phzvl_i[10][4]),
.phzvl_i_10_5_V(reg_phzvl_i[10][5]),
.phzvl_i_10_6_V(reg_phzvl_i[10][6]),
.phzvl_i_10_7_V(reg_phzvl_i[10][7]),
.phzvl_i_10_8_V(reg_phzvl_i[10][8]),
.phzvl_i_11_0_V(reg_phzvl_i[11][0]),
.phzvl_i_11_1_V(reg_phzvl_i[11][1]),
.phzvl_i_11_2_V(reg_phzvl_i[11][2]),
.phzvl_i_11_3_V(reg_phzvl_i[11][3]),
.phzvl_i_11_4_V(reg_phzvl_i[11][4]),
.phzvl_i_11_5_V(reg_phzvl_i[11][5]),
.phzvl_i_11_6_V(reg_phzvl_i[11][6]),
.phzvl_i_11_7_V(reg_phzvl_i[11][7]),
.phzvl_i_11_8_V(reg_phzvl_i[11][8]),
.phzvl_i_12_0_V(reg_phzvl_i[12][0]),
.phzvl_i_12_1_V(reg_phzvl_i[12][1]),
.phzvl_i_12_2_V(reg_phzvl_i[12][2]),
.phzvl_i_12_3_V(reg_phzvl_i[12][3]),
.phzvl_i_12_4_V(reg_phzvl_i[12][4]),
.phzvl_i_12_5_V(reg_phzvl_i[12][5]),
.phzvl_i_12_6_V(reg_phzvl_i[12][6]),
.phzvl_i_12_7_V(reg_phzvl_i[12][7]),
.phzvl_i_12_8_V(reg_phzvl_i[12][8]),
.ph_hit_i_0_0_V(reg_ph_hit_i[0][0]),
.ph_hit_i_0_1_V(reg_ph_hit_i[0][1]),
.ph_hit_i_0_2_V(reg_ph_hit_i[0][2]),
.ph_hit_i_0_3_V(reg_ph_hit_i[0][3]),
.ph_hit_i_0_4_V(reg_ph_hit_i[0][4]),
.ph_hit_i_0_5_V(reg_ph_hit_i[0][5]),
.ph_hit_i_0_6_V(reg_ph_hit_i[0][6]),
.ph_hit_i_0_7_V(reg_ph_hit_i[0][7]),
.ph_hit_i_0_8_V(reg_ph_hit_i[0][8]),
.ph_hit_i_1_0_V(reg_ph_hit_i[1][0]),
.ph_hit_i_1_1_V(reg_ph_hit_i[1][1]),
.ph_hit_i_1_2_V(reg_ph_hit_i[1][2]),
.ph_hit_i_1_3_V(reg_ph_hit_i[1][3]),
.ph_hit_i_1_4_V(reg_ph_hit_i[1][4]),
.ph_hit_i_1_5_V(reg_ph_hit_i[1][5]),
.ph_hit_i_1_6_V(reg_ph_hit_i[1][6]),
.ph_hit_i_1_7_V(reg_ph_hit_i[1][7]),
.ph_hit_i_1_8_V(reg_ph_hit_i[1][8]),
.ph_hit_i_2_0_V(reg_ph_hit_i[2][0]),
.ph_hit_i_2_1_V(reg_ph_hit_i[2][1]),
.ph_hit_i_2_2_V(reg_ph_hit_i[2][2]),
.ph_hit_i_2_3_V(reg_ph_hit_i[2][3]),
.ph_hit_i_2_4_V(reg_ph_hit_i[2][4]),
.ph_hit_i_2_5_V(reg_ph_hit_i[2][5]),
.ph_hit_i_2_6_V(reg_ph_hit_i[2][6]),
.ph_hit_i_2_7_V(reg_ph_hit_i[2][7]),
.ph_hit_i_2_8_V(reg_ph_hit_i[2][8]),
.ph_hit_i_3_0_V(reg_ph_hit_i[3][0]),
.ph_hit_i_3_1_V(reg_ph_hit_i[3][1]),
.ph_hit_i_3_2_V(reg_ph_hit_i[3][2]),
.ph_hit_i_3_3_V(reg_ph_hit_i[3][3]),
.ph_hit_i_3_4_V(reg_ph_hit_i[3][4]),
.ph_hit_i_3_5_V(reg_ph_hit_i[3][5]),
.ph_hit_i_3_6_V(reg_ph_hit_i[3][6]),
.ph_hit_i_3_7_V(reg_ph_hit_i[3][7]),
.ph_hit_i_3_8_V(reg_ph_hit_i[3][8]),
.ph_hit_i_4_0_V(reg_ph_hit_i[4][0]),
.ph_hit_i_4_1_V(reg_ph_hit_i[4][1]),
.ph_hit_i_4_2_V(reg_ph_hit_i[4][2]),
.ph_hit_i_4_3_V(reg_ph_hit_i[4][3]),
.ph_hit_i_4_4_V(reg_ph_hit_i[4][4]),
.ph_hit_i_4_5_V(reg_ph_hit_i[4][5]),
.ph_hit_i_4_6_V(reg_ph_hit_i[4][6]),
.ph_hit_i_4_7_V(reg_ph_hit_i[4][7]),
.ph_hit_i_4_8_V(reg_ph_hit_i[4][8]),
.ph_hit_i_5_0_V(reg_ph_hit_i[5][0]),
.ph_hit_i_5_1_V(reg_ph_hit_i[5][1]),
.ph_hit_i_5_2_V(reg_ph_hit_i[5][2]),
.ph_hit_i_5_3_V(reg_ph_hit_i[5][3]),
.ph_hit_i_5_4_V(reg_ph_hit_i[5][4]),
.ph_hit_i_5_5_V(reg_ph_hit_i[5][5]),
.ph_hit_i_5_6_V(reg_ph_hit_i[5][6]),
.ph_hit_i_5_7_V(reg_ph_hit_i[5][7]),
.ph_hit_i_5_8_V(reg_ph_hit_i[5][8]),
.ph_hit_i_6_0_V(reg_ph_hit_i[6][0]),
.ph_hit_i_6_1_V(reg_ph_hit_i[6][1]),
.ph_hit_i_6_2_V(reg_ph_hit_i[6][2]),
.ph_hit_i_6_3_V(reg_ph_hit_i[6][3]),
.ph_hit_i_6_4_V(reg_ph_hit_i[6][4]),
.ph_hit_i_6_5_V(reg_ph_hit_i[6][5]),
.ph_hit_i_6_6_V(reg_ph_hit_i[6][6]),
.ph_hit_i_6_7_V(reg_ph_hit_i[6][7]),
.ph_hit_i_6_8_V(reg_ph_hit_i[6][8]),
.ph_hit_i_7_0_V(reg_ph_hit_i[7][0]),
.ph_hit_i_7_1_V(reg_ph_hit_i[7][1]),
.ph_hit_i_7_2_V(reg_ph_hit_i[7][2]),
.ph_hit_i_7_3_V(reg_ph_hit_i[7][3]),
.ph_hit_i_7_4_V(reg_ph_hit_i[7][4]),
.ph_hit_i_7_5_V(reg_ph_hit_i[7][5]),
.ph_hit_i_7_6_V(reg_ph_hit_i[7][6]),
.ph_hit_i_7_7_V(reg_ph_hit_i[7][7]),
.ph_hit_i_7_8_V(reg_ph_hit_i[7][8]),
.ph_hit_i_8_0_V(reg_ph_hit_i[8][0]),
.ph_hit_i_8_1_V(reg_ph_hit_i[8][1]),
.ph_hit_i_8_2_V(reg_ph_hit_i[8][2]),
.ph_hit_i_8_3_V(reg_ph_hit_i[8][3]),
.ph_hit_i_8_4_V(reg_ph_hit_i[8][4]),
.ph_hit_i_8_5_V(reg_ph_hit_i[8][5]),
.ph_hit_i_8_6_V(reg_ph_hit_i[8][6]),
.ph_hit_i_8_7_V(reg_ph_hit_i[8][7]),
.ph_hit_i_8_8_V(reg_ph_hit_i[8][8]),
.ph_hit_i_9_0_V(reg_ph_hit_i[9][0]),
.ph_hit_i_9_1_V(reg_ph_hit_i[9][1]),
.ph_hit_i_9_2_V(reg_ph_hit_i[9][2]),
.ph_hit_i_9_3_V(reg_ph_hit_i[9][3]),
.ph_hit_i_9_4_V(reg_ph_hit_i[9][4]),
.ph_hit_i_9_5_V(reg_ph_hit_i[9][5]),
.ph_hit_i_9_6_V(reg_ph_hit_i[9][6]),
.ph_hit_i_9_7_V(reg_ph_hit_i[9][7]),
.ph_hit_i_9_8_V(reg_ph_hit_i[9][8]),
.ph_hit_i_10_0_V(reg_ph_hit_i[10][0]),
.ph_hit_i_10_1_V(reg_ph_hit_i[10][1]),
.ph_hit_i_10_2_V(reg_ph_hit_i[10][2]),
.ph_hit_i_10_3_V(reg_ph_hit_i[10][3]),
.ph_hit_i_10_4_V(reg_ph_hit_i[10][4]),
.ph_hit_i_10_5_V(reg_ph_hit_i[10][5]),
.ph_hit_i_10_6_V(reg_ph_hit_i[10][6]),
.ph_hit_i_10_7_V(reg_ph_hit_i[10][7]),
.ph_hit_i_10_8_V(reg_ph_hit_i[10][8]),
.ph_hit_i_11_0_V(reg_ph_hit_i[11][0]),
.ph_hit_i_11_1_V(reg_ph_hit_i[11][1]),
.ph_hit_i_11_2_V(reg_ph_hit_i[11][2]),
.ph_hit_i_11_3_V(reg_ph_hit_i[11][3]),
.ph_hit_i_11_4_V(reg_ph_hit_i[11][4]),
.ph_hit_i_11_5_V(reg_ph_hit_i[11][5]),
.ph_hit_i_11_6_V(reg_ph_hit_i[11][6]),
.ph_hit_i_11_7_V(reg_ph_hit_i[11][7]),
.ph_hit_i_11_8_V(reg_ph_hit_i[11][8]),
.ph_hit_i_12_0_V(reg_ph_hit_i[12][0]),
.ph_hit_i_12_1_V(reg_ph_hit_i[12][1]),
.ph_hit_i_12_2_V(reg_ph_hit_i[12][2]),
.ph_hit_i_12_3_V(reg_ph_hit_i[12][3]),
.ph_hit_i_12_4_V(reg_ph_hit_i[12][4]),
.ph_hit_i_12_5_V(reg_ph_hit_i[12][5]),
.ph_hit_i_12_6_V(reg_ph_hit_i[12][6]),
.ph_hit_i_12_7_V(reg_ph_hit_i[12][7]),
.ph_hit_i_12_8_V(reg_ph_hit_i[12][8]),
.time_o_0_0_0_0_V(wire_time_o[0][0][0][0]),
.time_o_0_0_0_1_V(wire_time_o[0][0][0][1]),
.time_o_0_0_1_0_V(wire_time_o[0][0][1][0]),
.time_o_0_0_1_1_V(wire_time_o[0][0][1][1]),
.time_o_0_0_2_0_V(wire_time_o[0][0][2][0]),
.time_o_0_0_2_1_V(wire_time_o[0][0][2][1]),
.time_o_0_0_3_0_V(wire_time_o[0][0][3][0]),
.time_o_0_0_3_1_V(wire_time_o[0][0][3][1]),
.time_o_0_0_4_0_V(wire_time_o[0][0][4][0]),
.time_o_0_0_4_1_V(wire_time_o[0][0][4][1]),
.time_o_0_0_5_0_V(wire_time_o[0][0][5][0]),
.time_o_0_0_5_1_V(wire_time_o[0][0][5][1]),
.time_o_0_0_6_0_V(wire_time_o[0][0][6][0]),
.time_o_0_0_6_1_V(wire_time_o[0][0][6][1]),
.time_o_0_0_7_0_V(wire_time_o[0][0][7][0]),
.time_o_0_0_7_1_V(wire_time_o[0][0][7][1]),
.time_o_0_0_8_0_V(wire_time_o[0][0][8][0]),
.time_o_0_0_8_1_V(wire_time_o[0][0][8][1]),
.time_o_0_1_0_0_V(wire_time_o[0][1][0][0]),
.time_o_0_1_0_1_V(wire_time_o[0][1][0][1]),
.time_o_0_1_1_0_V(wire_time_o[0][1][1][0]),
.time_o_0_1_1_1_V(wire_time_o[0][1][1][1]),
.time_o_0_1_2_0_V(wire_time_o[0][1][2][0]),
.time_o_0_1_2_1_V(wire_time_o[0][1][2][1]),
.time_o_0_1_3_0_V(wire_time_o[0][1][3][0]),
.time_o_0_1_3_1_V(wire_time_o[0][1][3][1]),
.time_o_0_1_4_0_V(wire_time_o[0][1][4][0]),
.time_o_0_1_4_1_V(wire_time_o[0][1][4][1]),
.time_o_0_1_5_0_V(wire_time_o[0][1][5][0]),
.time_o_0_1_5_1_V(wire_time_o[0][1][5][1]),
.time_o_0_1_6_0_V(wire_time_o[0][1][6][0]),
.time_o_0_1_6_1_V(wire_time_o[0][1][6][1]),
.time_o_0_1_7_0_V(wire_time_o[0][1][7][0]),
.time_o_0_1_7_1_V(wire_time_o[0][1][7][1]),
.time_o_0_1_8_0_V(wire_time_o[0][1][8][0]),
.time_o_0_1_8_1_V(wire_time_o[0][1][8][1]),
.time_o_0_2_0_0_V(wire_time_o[0][2][0][0]),
.time_o_0_2_0_1_V(wire_time_o[0][2][0][1]),
.time_o_0_2_1_0_V(wire_time_o[0][2][1][0]),
.time_o_0_2_1_1_V(wire_time_o[0][2][1][1]),
.time_o_0_2_2_0_V(wire_time_o[0][2][2][0]),
.time_o_0_2_2_1_V(wire_time_o[0][2][2][1]),
.time_o_0_2_3_0_V(wire_time_o[0][2][3][0]),
.time_o_0_2_3_1_V(wire_time_o[0][2][3][1]),
.time_o_0_2_4_0_V(wire_time_o[0][2][4][0]),
.time_o_0_2_4_1_V(wire_time_o[0][2][4][1]),
.time_o_0_2_5_0_V(wire_time_o[0][2][5][0]),
.time_o_0_2_5_1_V(wire_time_o[0][2][5][1]),
.time_o_0_2_6_0_V(wire_time_o[0][2][6][0]),
.time_o_0_2_6_1_V(wire_time_o[0][2][6][1]),
.time_o_0_2_7_0_V(wire_time_o[0][2][7][0]),
.time_o_0_2_7_1_V(wire_time_o[0][2][7][1]),
.time_o_0_2_8_0_V(wire_time_o[0][2][8][0]),
.time_o_0_2_8_1_V(wire_time_o[0][2][8][1]),
.time_o_0_3_0_0_V(wire_time_o[0][3][0][0]),
.time_o_0_3_0_1_V(wire_time_o[0][3][0][1]),
.time_o_0_3_1_0_V(wire_time_o[0][3][1][0]),
.time_o_0_3_1_1_V(wire_time_o[0][3][1][1]),
.time_o_0_3_2_0_V(wire_time_o[0][3][2][0]),
.time_o_0_3_2_1_V(wire_time_o[0][3][2][1]),
.time_o_0_3_3_0_V(wire_time_o[0][3][3][0]),
.time_o_0_3_3_1_V(wire_time_o[0][3][3][1]),
.time_o_0_3_4_0_V(wire_time_o[0][3][4][0]),
.time_o_0_3_4_1_V(wire_time_o[0][3][4][1]),
.time_o_0_3_5_0_V(wire_time_o[0][3][5][0]),
.time_o_0_3_5_1_V(wire_time_o[0][3][5][1]),
.time_o_0_3_6_0_V(wire_time_o[0][3][6][0]),
.time_o_0_3_6_1_V(wire_time_o[0][3][6][1]),
.time_o_0_3_7_0_V(wire_time_o[0][3][7][0]),
.time_o_0_3_7_1_V(wire_time_o[0][3][7][1]),
.time_o_0_3_8_0_V(wire_time_o[0][3][8][0]),
.time_o_0_3_8_1_V(wire_time_o[0][3][8][1]),
.time_o_0_4_0_0_V(wire_time_o[0][4][0][0]),
.time_o_0_4_0_1_V(wire_time_o[0][4][0][1]),
.time_o_0_4_1_0_V(wire_time_o[0][4][1][0]),
.time_o_0_4_1_1_V(wire_time_o[0][4][1][1]),
.time_o_0_4_2_0_V(wire_time_o[0][4][2][0]),
.time_o_0_4_2_1_V(wire_time_o[0][4][2][1]),
.time_o_0_4_3_0_V(wire_time_o[0][4][3][0]),
.time_o_0_4_3_1_V(wire_time_o[0][4][3][1]),
.time_o_0_4_4_0_V(wire_time_o[0][4][4][0]),
.time_o_0_4_4_1_V(wire_time_o[0][4][4][1]),
.time_o_0_4_5_0_V(wire_time_o[0][4][5][0]),
.time_o_0_4_5_1_V(wire_time_o[0][4][5][1]),
.time_o_0_4_6_0_V(wire_time_o[0][4][6][0]),
.time_o_0_4_6_1_V(wire_time_o[0][4][6][1]),
.time_o_0_4_7_0_V(wire_time_o[0][4][7][0]),
.time_o_0_4_7_1_V(wire_time_o[0][4][7][1]),
.time_o_0_4_8_0_V(wire_time_o[0][4][8][0]),
.time_o_0_4_8_1_V(wire_time_o[0][4][8][1]),
.time_o_0_5_0_0_V(wire_time_o[0][5][0][0]),
.time_o_0_5_0_1_V(wire_time_o[0][5][0][1]),
.time_o_0_5_1_0_V(wire_time_o[0][5][1][0]),
.time_o_0_5_1_1_V(wire_time_o[0][5][1][1]),
.time_o_0_5_2_0_V(wire_time_o[0][5][2][0]),
.time_o_0_5_2_1_V(wire_time_o[0][5][2][1]),
.time_o_0_5_3_0_V(wire_time_o[0][5][3][0]),
.time_o_0_5_3_1_V(wire_time_o[0][5][3][1]),
.time_o_0_5_4_0_V(wire_time_o[0][5][4][0]),
.time_o_0_5_4_1_V(wire_time_o[0][5][4][1]),
.time_o_0_5_5_0_V(wire_time_o[0][5][5][0]),
.time_o_0_5_5_1_V(wire_time_o[0][5][5][1]),
.time_o_0_5_6_0_V(wire_time_o[0][5][6][0]),
.time_o_0_5_6_1_V(wire_time_o[0][5][6][1]),
.time_o_0_5_7_0_V(wire_time_o[0][5][7][0]),
.time_o_0_5_7_1_V(wire_time_o[0][5][7][1]),
.time_o_0_5_8_0_V(wire_time_o[0][5][8][0]),
.time_o_0_5_8_1_V(wire_time_o[0][5][8][1]),
.time_o_0_6_0_0_V(wire_time_o[0][6][0][0]),
.time_o_0_6_0_1_V(wire_time_o[0][6][0][1]),
.time_o_0_6_1_0_V(wire_time_o[0][6][1][0]),
.time_o_0_6_1_1_V(wire_time_o[0][6][1][1]),
.time_o_0_6_2_0_V(wire_time_o[0][6][2][0]),
.time_o_0_6_2_1_V(wire_time_o[0][6][2][1]),
.time_o_0_6_3_0_V(wire_time_o[0][6][3][0]),
.time_o_0_6_3_1_V(wire_time_o[0][6][3][1]),
.time_o_0_6_4_0_V(wire_time_o[0][6][4][0]),
.time_o_0_6_4_1_V(wire_time_o[0][6][4][1]),
.time_o_0_6_5_0_V(wire_time_o[0][6][5][0]),
.time_o_0_6_5_1_V(wire_time_o[0][6][5][1]),
.time_o_0_6_6_0_V(wire_time_o[0][6][6][0]),
.time_o_0_6_6_1_V(wire_time_o[0][6][6][1]),
.time_o_0_6_7_0_V(wire_time_o[0][6][7][0]),
.time_o_0_6_7_1_V(wire_time_o[0][6][7][1]),
.time_o_0_6_8_0_V(wire_time_o[0][6][8][0]),
.time_o_0_6_8_1_V(wire_time_o[0][6][8][1]),
.vl_o_0_0_0_V(wire_vl_o[0][0][0]),
.vl_o_0_0_1_V(wire_vl_o[0][0][1]),
.vl_o_0_0_2_V(wire_vl_o[0][0][2]),
.vl_o_0_0_3_V(wire_vl_o[0][0][3]),
.vl_o_0_0_4_V(wire_vl_o[0][0][4]),
.vl_o_0_0_5_V(wire_vl_o[0][0][5]),
.vl_o_0_0_6_V(wire_vl_o[0][0][6]),
.vl_o_0_0_7_V(wire_vl_o[0][0][7]),
.vl_o_0_0_8_V(wire_vl_o[0][0][8]),
.vl_o_0_1_0_V(wire_vl_o[0][1][0]),
.vl_o_0_1_1_V(wire_vl_o[0][1][1]),
.vl_o_0_1_2_V(wire_vl_o[0][1][2]),
.vl_o_0_1_3_V(wire_vl_o[0][1][3]),
.vl_o_0_1_4_V(wire_vl_o[0][1][4]),
.vl_o_0_1_5_V(wire_vl_o[0][1][5]),
.vl_o_0_1_6_V(wire_vl_o[0][1][6]),
.vl_o_0_1_7_V(wire_vl_o[0][1][7]),
.vl_o_0_1_8_V(wire_vl_o[0][1][8]),
.vl_o_0_2_0_V(wire_vl_o[0][2][0]),
.vl_o_0_2_1_V(wire_vl_o[0][2][1]),
.vl_o_0_2_2_V(wire_vl_o[0][2][2]),
.vl_o_0_2_3_V(wire_vl_o[0][2][3]),
.vl_o_0_2_4_V(wire_vl_o[0][2][4]),
.vl_o_0_2_5_V(wire_vl_o[0][2][5]),
.vl_o_0_2_6_V(wire_vl_o[0][2][6]),
.vl_o_0_2_7_V(wire_vl_o[0][2][7]),
.vl_o_0_2_8_V(wire_vl_o[0][2][8]),
.vl_o_0_3_0_V(wire_vl_o[0][3][0]),
.vl_o_0_3_1_V(wire_vl_o[0][3][1]),
.vl_o_0_3_2_V(wire_vl_o[0][3][2]),
.vl_o_0_3_3_V(wire_vl_o[0][3][3]),
.vl_o_0_3_4_V(wire_vl_o[0][3][4]),
.vl_o_0_3_5_V(wire_vl_o[0][3][5]),
.vl_o_0_3_6_V(wire_vl_o[0][3][6]),
.vl_o_0_3_7_V(wire_vl_o[0][3][7]),
.vl_o_0_3_8_V(wire_vl_o[0][3][8]),
.vl_o_0_4_0_V(wire_vl_o[0][4][0]),
.vl_o_0_4_1_V(wire_vl_o[0][4][1]),
.vl_o_0_4_2_V(wire_vl_o[0][4][2]),
.vl_o_0_4_3_V(wire_vl_o[0][4][3]),
.vl_o_0_4_4_V(wire_vl_o[0][4][4]),
.vl_o_0_4_5_V(wire_vl_o[0][4][5]),
.vl_o_0_4_6_V(wire_vl_o[0][4][6]),
.vl_o_0_4_7_V(wire_vl_o[0][4][7]),
.vl_o_0_4_8_V(wire_vl_o[0][4][8]),
.vl_o_0_5_0_V(wire_vl_o[0][5][0]),
.vl_o_0_5_1_V(wire_vl_o[0][5][1]),
.vl_o_0_5_2_V(wire_vl_o[0][5][2]),
.vl_o_0_5_3_V(wire_vl_o[0][5][3]),
.vl_o_0_5_4_V(wire_vl_o[0][5][4]),
.vl_o_0_5_5_V(wire_vl_o[0][5][5]),
.vl_o_0_5_6_V(wire_vl_o[0][5][6]),
.vl_o_0_5_7_V(wire_vl_o[0][5][7]),
.vl_o_0_5_8_V(wire_vl_o[0][5][8]),
.vl_o_0_6_0_V(wire_vl_o[0][6][0]),
.vl_o_0_6_1_V(wire_vl_o[0][6][1]),
.vl_o_0_6_2_V(wire_vl_o[0][6][2]),
.vl_o_0_6_3_V(wire_vl_o[0][6][3]),
.vl_o_0_6_4_V(wire_vl_o[0][6][4]),
.vl_o_0_6_5_V(wire_vl_o[0][6][5]),
.vl_o_0_6_6_V(wire_vl_o[0][6][6]),
.vl_o_0_6_7_V(wire_vl_o[0][6][7]),
.vl_o_0_6_8_V(wire_vl_o[0][6][8]),
.vl_o_0_7_0_V(wire_vl_o[0][7][0]),
.vl_o_0_7_1_V(wire_vl_o[0][7][1]),
.vl_o_0_7_2_V(wire_vl_o[0][7][2]),
.vl_o_0_7_3_V(wire_vl_o[0][7][3]),
.vl_o_0_7_4_V(wire_vl_o[0][7][4]),
.vl_o_0_7_5_V(wire_vl_o[0][7][5]),
.vl_o_0_7_6_V(wire_vl_o[0][7][6]),
.vl_o_0_7_7_V(wire_vl_o[0][7][7]),
.vl_o_0_7_8_V(wire_vl_o[0][7][8]),
.vl_o_0_8_0_V(wire_vl_o[0][8][0]),
.vl_o_0_8_1_V(wire_vl_o[0][8][1]),
.vl_o_0_8_2_V(wire_vl_o[0][8][2]),
.vl_o_0_8_3_V(wire_vl_o[0][8][3]),
.vl_o_0_8_4_V(wire_vl_o[0][8][4]),
.vl_o_0_8_5_V(wire_vl_o[0][8][5]),
.vl_o_0_8_6_V(wire_vl_o[0][8][6]),
.vl_o_0_8_7_V(wire_vl_o[0][8][7]),
.vl_o_0_8_8_V(wire_vl_o[0][8][8]),
.vl_o_0_9_0_V(wire_vl_o[0][9][0]),
.vl_o_0_9_1_V(wire_vl_o[0][9][1]),
.vl_o_0_9_2_V(wire_vl_o[0][9][2]),
.vl_o_0_9_3_V(wire_vl_o[0][9][3]),
.vl_o_0_9_4_V(wire_vl_o[0][9][4]),
.vl_o_0_9_5_V(wire_vl_o[0][9][5]),
.vl_o_0_9_6_V(wire_vl_o[0][9][6]),
.vl_o_0_9_7_V(wire_vl_o[0][9][7]),
.vl_o_0_9_8_V(wire_vl_o[0][9][8]),
.vl_o_0_10_0_V(wire_vl_o[0][10][0]),
.vl_o_0_10_1_V(wire_vl_o[0][10][1]),
.vl_o_0_10_2_V(wire_vl_o[0][10][2]),
.vl_o_0_10_3_V(wire_vl_o[0][10][3]),
.vl_o_0_10_4_V(wire_vl_o[0][10][4]),
.vl_o_0_10_5_V(wire_vl_o[0][10][5]),
.vl_o_0_10_6_V(wire_vl_o[0][10][6]),
.vl_o_0_10_7_V(wire_vl_o[0][10][7]),
.vl_o_0_10_8_V(wire_vl_o[0][10][8]),
.vl_o_0_11_0_V(wire_vl_o[0][11][0]),
.vl_o_0_11_1_V(wire_vl_o[0][11][1]),
.vl_o_0_11_2_V(wire_vl_o[0][11][2]),
.vl_o_0_11_3_V(wire_vl_o[0][11][3]),
.vl_o_0_11_4_V(wire_vl_o[0][11][4]),
.vl_o_0_11_5_V(wire_vl_o[0][11][5]),
.vl_o_0_11_6_V(wire_vl_o[0][11][6]),
.vl_o_0_11_7_V(wire_vl_o[0][11][7]),
.vl_o_0_11_8_V(wire_vl_o[0][11][8]),
.vl_o_0_12_0_V(wire_vl_o[0][12][0]),
.vl_o_0_12_1_V(wire_vl_o[0][12][1]),
.vl_o_0_12_2_V(wire_vl_o[0][12][2]),
.vl_o_0_12_3_V(wire_vl_o[0][12][3]),
.vl_o_0_12_4_V(wire_vl_o[0][12][4]),
.vl_o_0_12_5_V(wire_vl_o[0][12][5]),
.vl_o_0_12_6_V(wire_vl_o[0][12][6]),
.vl_o_0_12_7_V(wire_vl_o[0][12][7]),
.vl_o_0_12_8_V(wire_vl_o[0][12][8]),
.q_o_0_0_0_0_V(wire_q_o[0][0][0][0]),
.q_o_0_0_0_1_V(wire_q_o[0][0][0][1]),
.q_o_0_0_0_2_V(wire_q_o[0][0][0][2]),
.q_o_0_0_1_0_V(wire_q_o[0][0][1][0]),
.q_o_0_0_1_1_V(wire_q_o[0][0][1][1]),
.q_o_0_0_1_2_V(wire_q_o[0][0][1][2]),
.q_o_0_0_2_0_V(wire_q_o[0][0][2][0]),
.q_o_0_0_2_1_V(wire_q_o[0][0][2][1]),
.q_o_0_0_2_2_V(wire_q_o[0][0][2][2]),
.q_o_0_0_3_0_V(wire_q_o[0][0][3][0]),
.q_o_0_0_3_1_V(wire_q_o[0][0][3][1]),
.q_o_0_0_3_2_V(wire_q_o[0][0][3][2]),
.q_o_0_0_4_0_V(wire_q_o[0][0][4][0]),
.q_o_0_0_4_1_V(wire_q_o[0][0][4][1]),
.q_o_0_0_4_2_V(wire_q_o[0][0][4][2]),
.q_o_0_0_5_0_V(wire_q_o[0][0][5][0]),
.q_o_0_0_5_1_V(wire_q_o[0][0][5][1]),
.q_o_0_0_5_2_V(wire_q_o[0][0][5][2]),
.q_o_0_0_6_0_V(wire_q_o[0][0][6][0]),
.q_o_0_0_6_1_V(wire_q_o[0][0][6][1]),
.q_o_0_0_6_2_V(wire_q_o[0][0][6][2]),
.q_o_0_0_7_0_V(wire_q_o[0][0][7][0]),
.q_o_0_0_7_1_V(wire_q_o[0][0][7][1]),
.q_o_0_0_7_2_V(wire_q_o[0][0][7][2]),
.q_o_0_0_8_0_V(wire_q_o[0][0][8][0]),
.q_o_0_0_8_1_V(wire_q_o[0][0][8][1]),
.q_o_0_0_8_2_V(wire_q_o[0][0][8][2]),
.q_o_0_1_0_0_V(wire_q_o[0][1][0][0]),
.q_o_0_1_0_1_V(wire_q_o[0][1][0][1]),
.q_o_0_1_0_2_V(wire_q_o[0][1][0][2]),
.q_o_0_1_1_0_V(wire_q_o[0][1][1][0]),
.q_o_0_1_1_1_V(wire_q_o[0][1][1][1]),
.q_o_0_1_1_2_V(wire_q_o[0][1][1][2]),
.q_o_0_1_2_0_V(wire_q_o[0][1][2][0]),
.q_o_0_1_2_1_V(wire_q_o[0][1][2][1]),
.q_o_0_1_2_2_V(wire_q_o[0][1][2][2]),
.q_o_0_1_3_0_V(wire_q_o[0][1][3][0]),
.q_o_0_1_3_1_V(wire_q_o[0][1][3][1]),
.q_o_0_1_3_2_V(wire_q_o[0][1][3][2]),
.q_o_0_1_4_0_V(wire_q_o[0][1][4][0]),
.q_o_0_1_4_1_V(wire_q_o[0][1][4][1]),
.q_o_0_1_4_2_V(wire_q_o[0][1][4][2]),
.q_o_0_1_5_0_V(wire_q_o[0][1][5][0]),
.q_o_0_1_5_1_V(wire_q_o[0][1][5][1]),
.q_o_0_1_5_2_V(wire_q_o[0][1][5][2]),
.q_o_0_1_6_0_V(wire_q_o[0][1][6][0]),
.q_o_0_1_6_1_V(wire_q_o[0][1][6][1]),
.q_o_0_1_6_2_V(wire_q_o[0][1][6][2]),
.q_o_0_1_7_0_V(wire_q_o[0][1][7][0]),
.q_o_0_1_7_1_V(wire_q_o[0][1][7][1]),
.q_o_0_1_7_2_V(wire_q_o[0][1][7][2]),
.q_o_0_1_8_0_V(wire_q_o[0][1][8][0]),
.q_o_0_1_8_1_V(wire_q_o[0][1][8][1]),
.q_o_0_1_8_2_V(wire_q_o[0][1][8][2]),
.q_o_0_2_0_0_V(wire_q_o[0][2][0][0]),
.q_o_0_2_0_1_V(wire_q_o[0][2][0][1]),
.q_o_0_2_0_2_V(wire_q_o[0][2][0][2]),
.q_o_0_2_1_0_V(wire_q_o[0][2][1][0]),
.q_o_0_2_1_1_V(wire_q_o[0][2][1][1]),
.q_o_0_2_1_2_V(wire_q_o[0][2][1][2]),
.q_o_0_2_2_0_V(wire_q_o[0][2][2][0]),
.q_o_0_2_2_1_V(wire_q_o[0][2][2][1]),
.q_o_0_2_2_2_V(wire_q_o[0][2][2][2]),
.q_o_0_2_3_0_V(wire_q_o[0][2][3][0]),
.q_o_0_2_3_1_V(wire_q_o[0][2][3][1]),
.q_o_0_2_3_2_V(wire_q_o[0][2][3][2]),
.q_o_0_2_4_0_V(wire_q_o[0][2][4][0]),
.q_o_0_2_4_1_V(wire_q_o[0][2][4][1]),
.q_o_0_2_4_2_V(wire_q_o[0][2][4][2]),
.q_o_0_2_5_0_V(wire_q_o[0][2][5][0]),
.q_o_0_2_5_1_V(wire_q_o[0][2][5][1]),
.q_o_0_2_5_2_V(wire_q_o[0][2][5][2]),
.q_o_0_2_6_0_V(wire_q_o[0][2][6][0]),
.q_o_0_2_6_1_V(wire_q_o[0][2][6][1]),
.q_o_0_2_6_2_V(wire_q_o[0][2][6][2]),
.q_o_0_2_7_0_V(wire_q_o[0][2][7][0]),
.q_o_0_2_7_1_V(wire_q_o[0][2][7][1]),
.q_o_0_2_7_2_V(wire_q_o[0][2][7][2]),
.q_o_0_2_8_0_V(wire_q_o[0][2][8][0]),
.q_o_0_2_8_1_V(wire_q_o[0][2][8][1]),
.q_o_0_2_8_2_V(wire_q_o[0][2][8][2]),
.q_o_0_3_0_0_V(wire_q_o[0][3][0][0]),
.q_o_0_3_0_1_V(wire_q_o[0][3][0][1]),
.q_o_0_3_0_2_V(wire_q_o[0][3][0][2]),
.q_o_0_3_1_0_V(wire_q_o[0][3][1][0]),
.q_o_0_3_1_1_V(wire_q_o[0][3][1][1]),
.q_o_0_3_1_2_V(wire_q_o[0][3][1][2]),
.q_o_0_3_2_0_V(wire_q_o[0][3][2][0]),
.q_o_0_3_2_1_V(wire_q_o[0][3][2][1]),
.q_o_0_3_2_2_V(wire_q_o[0][3][2][2]),
.q_o_0_3_3_0_V(wire_q_o[0][3][3][0]),
.q_o_0_3_3_1_V(wire_q_o[0][3][3][1]),
.q_o_0_3_3_2_V(wire_q_o[0][3][3][2]),
.q_o_0_3_4_0_V(wire_q_o[0][3][4][0]),
.q_o_0_3_4_1_V(wire_q_o[0][3][4][1]),
.q_o_0_3_4_2_V(wire_q_o[0][3][4][2]),
.q_o_0_3_5_0_V(wire_q_o[0][3][5][0]),
.q_o_0_3_5_1_V(wire_q_o[0][3][5][1]),
.q_o_0_3_5_2_V(wire_q_o[0][3][5][2]),
.q_o_0_3_6_0_V(wire_q_o[0][3][6][0]),
.q_o_0_3_6_1_V(wire_q_o[0][3][6][1]),
.q_o_0_3_6_2_V(wire_q_o[0][3][6][2]),
.q_o_0_3_7_0_V(wire_q_o[0][3][7][0]),
.q_o_0_3_7_1_V(wire_q_o[0][3][7][1]),
.q_o_0_3_7_2_V(wire_q_o[0][3][7][2]),
.q_o_0_3_8_0_V(wire_q_o[0][3][8][0]),
.q_o_0_3_8_1_V(wire_q_o[0][3][8][1]),
.q_o_0_3_8_2_V(wire_q_o[0][3][8][2]),
.q_o_0_4_0_0_V(wire_q_o[0][4][0][0]),
.q_o_0_4_0_1_V(wire_q_o[0][4][0][1]),
.q_o_0_4_0_2_V(wire_q_o[0][4][0][2]),
.q_o_0_4_1_0_V(wire_q_o[0][4][1][0]),
.q_o_0_4_1_1_V(wire_q_o[0][4][1][1]),
.q_o_0_4_1_2_V(wire_q_o[0][4][1][2]),
.q_o_0_4_2_0_V(wire_q_o[0][4][2][0]),
.q_o_0_4_2_1_V(wire_q_o[0][4][2][1]),
.q_o_0_4_2_2_V(wire_q_o[0][4][2][2]),
.q_o_0_4_3_0_V(wire_q_o[0][4][3][0]),
.q_o_0_4_3_1_V(wire_q_o[0][4][3][1]),
.q_o_0_4_3_2_V(wire_q_o[0][4][3][2]),
.q_o_0_4_4_0_V(wire_q_o[0][4][4][0]),
.q_o_0_4_4_1_V(wire_q_o[0][4][4][1]),
.q_o_0_4_4_2_V(wire_q_o[0][4][4][2]),
.q_o_0_4_5_0_V(wire_q_o[0][4][5][0]),
.q_o_0_4_5_1_V(wire_q_o[0][4][5][1]),
.q_o_0_4_5_2_V(wire_q_o[0][4][5][2]),
.q_o_0_4_6_0_V(wire_q_o[0][4][6][0]),
.q_o_0_4_6_1_V(wire_q_o[0][4][6][1]),
.q_o_0_4_6_2_V(wire_q_o[0][4][6][2]),
.q_o_0_4_7_0_V(wire_q_o[0][4][7][0]),
.q_o_0_4_7_1_V(wire_q_o[0][4][7][1]),
.q_o_0_4_7_2_V(wire_q_o[0][4][7][2]),
.q_o_0_4_8_0_V(wire_q_o[0][4][8][0]),
.q_o_0_4_8_1_V(wire_q_o[0][4][8][1]),
.q_o_0_4_8_2_V(wire_q_o[0][4][8][2]),
.q_o_0_5_0_0_V(wire_q_o[0][5][0][0]),
.q_o_0_5_0_1_V(wire_q_o[0][5][0][1]),
.q_o_0_5_0_2_V(wire_q_o[0][5][0][2]),
.q_o_0_5_1_0_V(wire_q_o[0][5][1][0]),
.q_o_0_5_1_1_V(wire_q_o[0][5][1][1]),
.q_o_0_5_1_2_V(wire_q_o[0][5][1][2]),
.q_o_0_5_2_0_V(wire_q_o[0][5][2][0]),
.q_o_0_5_2_1_V(wire_q_o[0][5][2][1]),
.q_o_0_5_2_2_V(wire_q_o[0][5][2][2]),
.q_o_0_5_3_0_V(wire_q_o[0][5][3][0]),
.q_o_0_5_3_1_V(wire_q_o[0][5][3][1]),
.q_o_0_5_3_2_V(wire_q_o[0][5][3][2]),
.q_o_0_5_4_0_V(wire_q_o[0][5][4][0]),
.q_o_0_5_4_1_V(wire_q_o[0][5][4][1]),
.q_o_0_5_4_2_V(wire_q_o[0][5][4][2]),
.q_o_0_5_5_0_V(wire_q_o[0][5][5][0]),
.q_o_0_5_5_1_V(wire_q_o[0][5][5][1]),
.q_o_0_5_5_2_V(wire_q_o[0][5][5][2]),
.q_o_0_5_6_0_V(wire_q_o[0][5][6][0]),
.q_o_0_5_6_1_V(wire_q_o[0][5][6][1]),
.q_o_0_5_6_2_V(wire_q_o[0][5][6][2]),
.q_o_0_5_7_0_V(wire_q_o[0][5][7][0]),
.q_o_0_5_7_1_V(wire_q_o[0][5][7][1]),
.q_o_0_5_7_2_V(wire_q_o[0][5][7][2]),
.q_o_0_5_8_0_V(wire_q_o[0][5][8][0]),
.q_o_0_5_8_1_V(wire_q_o[0][5][8][1]),
.q_o_0_5_8_2_V(wire_q_o[0][5][8][2]),
.q_o_0_6_0_0_V(wire_q_o[0][6][0][0]),
.q_o_0_6_0_1_V(wire_q_o[0][6][0][1]),
.q_o_0_6_0_2_V(wire_q_o[0][6][0][2]),
.q_o_0_6_1_0_V(wire_q_o[0][6][1][0]),
.q_o_0_6_1_1_V(wire_q_o[0][6][1][1]),
.q_o_0_6_1_2_V(wire_q_o[0][6][1][2]),
.q_o_0_6_2_0_V(wire_q_o[0][6][2][0]),
.q_o_0_6_2_1_V(wire_q_o[0][6][2][1]),
.q_o_0_6_2_2_V(wire_q_o[0][6][2][2]),
.q_o_0_6_3_0_V(wire_q_o[0][6][3][0]),
.q_o_0_6_3_1_V(wire_q_o[0][6][3][1]),
.q_o_0_6_3_2_V(wire_q_o[0][6][3][2]),
.q_o_0_6_4_0_V(wire_q_o[0][6][4][0]),
.q_o_0_6_4_1_V(wire_q_o[0][6][4][1]),
.q_o_0_6_4_2_V(wire_q_o[0][6][4][2]),
.q_o_0_6_5_0_V(wire_q_o[0][6][5][0]),
.q_o_0_6_5_1_V(wire_q_o[0][6][5][1]),
.q_o_0_6_5_2_V(wire_q_o[0][6][5][2]),
.q_o_0_6_6_0_V(wire_q_o[0][6][6][0]),
.q_o_0_6_6_1_V(wire_q_o[0][6][6][1]),
.q_o_0_6_6_2_V(wire_q_o[0][6][6][2]),
.q_o_0_6_7_0_V(wire_q_o[0][6][7][0]),
.q_o_0_6_7_1_V(wire_q_o[0][6][7][1]),
.q_o_0_6_7_2_V(wire_q_o[0][6][7][2]),
.q_o_0_6_8_0_V(wire_q_o[0][6][8][0]),
.q_o_0_6_8_1_V(wire_q_o[0][6][8][1]),
.q_o_0_6_8_2_V(wire_q_o[0][6][8][2]),
.q_o_0_7_0_0_V(wire_q_o[0][7][0][0]),
.q_o_0_7_0_1_V(wire_q_o[0][7][0][1]),
.q_o_0_7_0_2_V(wire_q_o[0][7][0][2]),
.q_o_0_7_1_0_V(wire_q_o[0][7][1][0]),
.q_o_0_7_1_1_V(wire_q_o[0][7][1][1]),
.q_o_0_7_1_2_V(wire_q_o[0][7][1][2]),
.q_o_0_7_2_0_V(wire_q_o[0][7][2][0]),
.q_o_0_7_2_1_V(wire_q_o[0][7][2][1]),
.q_o_0_7_2_2_V(wire_q_o[0][7][2][2]),
.q_o_0_7_3_0_V(wire_q_o[0][7][3][0]),
.q_o_0_7_3_1_V(wire_q_o[0][7][3][1]),
.q_o_0_7_3_2_V(wire_q_o[0][7][3][2]),
.q_o_0_7_4_0_V(wire_q_o[0][7][4][0]),
.q_o_0_7_4_1_V(wire_q_o[0][7][4][1]),
.q_o_0_7_4_2_V(wire_q_o[0][7][4][2]),
.q_o_0_7_5_0_V(wire_q_o[0][7][5][0]),
.q_o_0_7_5_1_V(wire_q_o[0][7][5][1]),
.q_o_0_7_5_2_V(wire_q_o[0][7][5][2]),
.q_o_0_7_6_0_V(wire_q_o[0][7][6][0]),
.q_o_0_7_6_1_V(wire_q_o[0][7][6][1]),
.q_o_0_7_6_2_V(wire_q_o[0][7][6][2]),
.q_o_0_7_7_0_V(wire_q_o[0][7][7][0]),
.q_o_0_7_7_1_V(wire_q_o[0][7][7][1]),
.q_o_0_7_7_2_V(wire_q_o[0][7][7][2]),
.q_o_0_7_8_0_V(wire_q_o[0][7][8][0]),
.q_o_0_7_8_1_V(wire_q_o[0][7][8][1]),
.q_o_0_7_8_2_V(wire_q_o[0][7][8][2]),
.q_o_0_8_0_0_V(wire_q_o[0][8][0][0]),
.q_o_0_8_0_1_V(wire_q_o[0][8][0][1]),
.q_o_0_8_0_2_V(wire_q_o[0][8][0][2]),
.q_o_0_8_1_0_V(wire_q_o[0][8][1][0]),
.q_o_0_8_1_1_V(wire_q_o[0][8][1][1]),
.q_o_0_8_1_2_V(wire_q_o[0][8][1][2]),
.q_o_0_8_2_0_V(wire_q_o[0][8][2][0]),
.q_o_0_8_2_1_V(wire_q_o[0][8][2][1]),
.q_o_0_8_2_2_V(wire_q_o[0][8][2][2]),
.q_o_0_8_3_0_V(wire_q_o[0][8][3][0]),
.q_o_0_8_3_1_V(wire_q_o[0][8][3][1]),
.q_o_0_8_3_2_V(wire_q_o[0][8][3][2]),
.q_o_0_8_4_0_V(wire_q_o[0][8][4][0]),
.q_o_0_8_4_1_V(wire_q_o[0][8][4][1]),
.q_o_0_8_4_2_V(wire_q_o[0][8][4][2]),
.q_o_0_8_5_0_V(wire_q_o[0][8][5][0]),
.q_o_0_8_5_1_V(wire_q_o[0][8][5][1]),
.q_o_0_8_5_2_V(wire_q_o[0][8][5][2]),
.q_o_0_8_6_0_V(wire_q_o[0][8][6][0]),
.q_o_0_8_6_1_V(wire_q_o[0][8][6][1]),
.q_o_0_8_6_2_V(wire_q_o[0][8][6][2]),
.q_o_0_8_7_0_V(wire_q_o[0][8][7][0]),
.q_o_0_8_7_1_V(wire_q_o[0][8][7][1]),
.q_o_0_8_7_2_V(wire_q_o[0][8][7][2]),
.q_o_0_8_8_0_V(wire_q_o[0][8][8][0]),
.q_o_0_8_8_1_V(wire_q_o[0][8][8][1]),
.q_o_0_8_8_2_V(wire_q_o[0][8][8][2]),
.q_o_0_9_0_0_V(wire_q_o[0][9][0][0]),
.q_o_0_9_0_1_V(wire_q_o[0][9][0][1]),
.q_o_0_9_0_2_V(wire_q_o[0][9][0][2]),
.q_o_0_9_1_0_V(wire_q_o[0][9][1][0]),
.q_o_0_9_1_1_V(wire_q_o[0][9][1][1]),
.q_o_0_9_1_2_V(wire_q_o[0][9][1][2]),
.q_o_0_9_2_0_V(wire_q_o[0][9][2][0]),
.q_o_0_9_2_1_V(wire_q_o[0][9][2][1]),
.q_o_0_9_2_2_V(wire_q_o[0][9][2][2]),
.q_o_0_9_3_0_V(wire_q_o[0][9][3][0]),
.q_o_0_9_3_1_V(wire_q_o[0][9][3][1]),
.q_o_0_9_3_2_V(wire_q_o[0][9][3][2]),
.q_o_0_9_4_0_V(wire_q_o[0][9][4][0]),
.q_o_0_9_4_1_V(wire_q_o[0][9][4][1]),
.q_o_0_9_4_2_V(wire_q_o[0][9][4][2]),
.q_o_0_9_5_0_V(wire_q_o[0][9][5][0]),
.q_o_0_9_5_1_V(wire_q_o[0][9][5][1]),
.q_o_0_9_5_2_V(wire_q_o[0][9][5][2]),
.q_o_0_9_6_0_V(wire_q_o[0][9][6][0]),
.q_o_0_9_6_1_V(wire_q_o[0][9][6][1]),
.q_o_0_9_6_2_V(wire_q_o[0][9][6][2]),
.q_o_0_9_7_0_V(wire_q_o[0][9][7][0]),
.q_o_0_9_7_1_V(wire_q_o[0][9][7][1]),
.q_o_0_9_7_2_V(wire_q_o[0][9][7][2]),
.q_o_0_9_8_0_V(wire_q_o[0][9][8][0]),
.q_o_0_9_8_1_V(wire_q_o[0][9][8][1]),
.q_o_0_9_8_2_V(wire_q_o[0][9][8][2]),
.q_o_0_10_0_0_V(wire_q_o[0][10][0][0]),
.q_o_0_10_0_1_V(wire_q_o[0][10][0][1]),
.q_o_0_10_0_2_V(wire_q_o[0][10][0][2]),
.q_o_0_10_1_0_V(wire_q_o[0][10][1][0]),
.q_o_0_10_1_1_V(wire_q_o[0][10][1][1]),
.q_o_0_10_1_2_V(wire_q_o[0][10][1][2]),
.q_o_0_10_2_0_V(wire_q_o[0][10][2][0]),
.q_o_0_10_2_1_V(wire_q_o[0][10][2][1]),
.q_o_0_10_2_2_V(wire_q_o[0][10][2][2]),
.q_o_0_10_3_0_V(wire_q_o[0][10][3][0]),
.q_o_0_10_3_1_V(wire_q_o[0][10][3][1]),
.q_o_0_10_3_2_V(wire_q_o[0][10][3][2]),
.q_o_0_10_4_0_V(wire_q_o[0][10][4][0]),
.q_o_0_10_4_1_V(wire_q_o[0][10][4][1]),
.q_o_0_10_4_2_V(wire_q_o[0][10][4][2]),
.q_o_0_10_5_0_V(wire_q_o[0][10][5][0]),
.q_o_0_10_5_1_V(wire_q_o[0][10][5][1]),
.q_o_0_10_5_2_V(wire_q_o[0][10][5][2]),
.q_o_0_10_6_0_V(wire_q_o[0][10][6][0]),
.q_o_0_10_6_1_V(wire_q_o[0][10][6][1]),
.q_o_0_10_6_2_V(wire_q_o[0][10][6][2]),
.q_o_0_10_7_0_V(wire_q_o[0][10][7][0]),
.q_o_0_10_7_1_V(wire_q_o[0][10][7][1]),
.q_o_0_10_7_2_V(wire_q_o[0][10][7][2]),
.q_o_0_10_8_0_V(wire_q_o[0][10][8][0]),
.q_o_0_10_8_1_V(wire_q_o[0][10][8][1]),
.q_o_0_10_8_2_V(wire_q_o[0][10][8][2]),
.q_o_0_11_0_0_V(wire_q_o[0][11][0][0]),
.q_o_0_11_0_1_V(wire_q_o[0][11][0][1]),
.q_o_0_11_0_2_V(wire_q_o[0][11][0][2]),
.q_o_0_11_1_0_V(wire_q_o[0][11][1][0]),
.q_o_0_11_1_1_V(wire_q_o[0][11][1][1]),
.q_o_0_11_1_2_V(wire_q_o[0][11][1][2]),
.q_o_0_11_2_0_V(wire_q_o[0][11][2][0]),
.q_o_0_11_2_1_V(wire_q_o[0][11][2][1]),
.q_o_0_11_2_2_V(wire_q_o[0][11][2][2]),
.q_o_0_11_3_0_V(wire_q_o[0][11][3][0]),
.q_o_0_11_3_1_V(wire_q_o[0][11][3][1]),
.q_o_0_11_3_2_V(wire_q_o[0][11][3][2]),
.q_o_0_11_4_0_V(wire_q_o[0][11][4][0]),
.q_o_0_11_4_1_V(wire_q_o[0][11][4][1]),
.q_o_0_11_4_2_V(wire_q_o[0][11][4][2]),
.q_o_0_11_5_0_V(wire_q_o[0][11][5][0]),
.q_o_0_11_5_1_V(wire_q_o[0][11][5][1]),
.q_o_0_11_5_2_V(wire_q_o[0][11][5][2]),
.q_o_0_11_6_0_V(wire_q_o[0][11][6][0]),
.q_o_0_11_6_1_V(wire_q_o[0][11][6][1]),
.q_o_0_11_6_2_V(wire_q_o[0][11][6][2]),
.q_o_0_11_7_0_V(wire_q_o[0][11][7][0]),
.q_o_0_11_7_1_V(wire_q_o[0][11][7][1]),
.q_o_0_11_7_2_V(wire_q_o[0][11][7][2]),
.q_o_0_11_8_0_V(wire_q_o[0][11][8][0]),
.q_o_0_11_8_1_V(wire_q_o[0][11][8][1]),
.q_o_0_11_8_2_V(wire_q_o[0][11][8][2]),
.q_o_0_12_0_0_V(wire_q_o[0][12][0][0]),
.q_o_0_12_0_1_V(wire_q_o[0][12][0][1]),
.q_o_0_12_0_2_V(wire_q_o[0][12][0][2]),
.q_o_0_12_1_0_V(wire_q_o[0][12][1][0]),
.q_o_0_12_1_1_V(wire_q_o[0][12][1][1]),
.q_o_0_12_1_2_V(wire_q_o[0][12][1][2]),
.q_o_0_12_2_0_V(wire_q_o[0][12][2][0]),
.q_o_0_12_2_1_V(wire_q_o[0][12][2][1]),
.q_o_0_12_2_2_V(wire_q_o[0][12][2][2]),
.q_o_0_12_3_0_V(wire_q_o[0][12][3][0]),
.q_o_0_12_3_1_V(wire_q_o[0][12][3][1]),
.q_o_0_12_3_2_V(wire_q_o[0][12][3][2]),
.q_o_0_12_4_0_V(wire_q_o[0][12][4][0]),
.q_o_0_12_4_1_V(wire_q_o[0][12][4][1]),
.q_o_0_12_4_2_V(wire_q_o[0][12][4][2]),
.q_o_0_12_5_0_V(wire_q_o[0][12][5][0]),
.q_o_0_12_5_1_V(wire_q_o[0][12][5][1]),
.q_o_0_12_5_2_V(wire_q_o[0][12][5][2]),
.q_o_0_12_6_0_V(wire_q_o[0][12][6][0]),
.q_o_0_12_6_1_V(wire_q_o[0][12][6][1]),
.q_o_0_12_6_2_V(wire_q_o[0][12][6][2]),
.q_o_0_12_7_0_V(wire_q_o[0][12][7][0]),
.q_o_0_12_7_1_V(wire_q_o[0][12][7][1]),
.q_o_0_12_7_2_V(wire_q_o[0][12][7][2]),
.q_o_0_12_8_0_V(wire_q_o[0][12][8][0]),
.q_o_0_12_8_1_V(wire_q_o[0][12][8][1]),
.q_o_0_12_8_2_V(wire_q_o[0][12][8][2]),
.cpatr_o_0_0_0_0_V(wire_cpatr_o[0][0][0][0]),
.cpatr_o_0_0_0_1_V(wire_cpatr_o[0][0][0][1]),
.cpatr_o_0_0_1_0_V(wire_cpatr_o[0][0][1][0]),
.cpatr_o_0_0_1_1_V(wire_cpatr_o[0][0][1][1]),
.cpatr_o_0_0_2_0_V(wire_cpatr_o[0][0][2][0]),
.cpatr_o_0_0_2_1_V(wire_cpatr_o[0][0][2][1]),
.cpatr_o_0_0_3_0_V(wire_cpatr_o[0][0][3][0]),
.cpatr_o_0_0_3_1_V(wire_cpatr_o[0][0][3][1]),
.cpatr_o_0_0_4_0_V(wire_cpatr_o[0][0][4][0]),
.cpatr_o_0_0_4_1_V(wire_cpatr_o[0][0][4][1]),
.cpatr_o_0_0_5_0_V(wire_cpatr_o[0][0][5][0]),
.cpatr_o_0_0_5_1_V(wire_cpatr_o[0][0][5][1]),
.cpatr_o_0_0_6_0_V(wire_cpatr_o[0][0][6][0]),
.cpatr_o_0_0_6_1_V(wire_cpatr_o[0][0][6][1]),
.cpatr_o_0_0_7_0_V(wire_cpatr_o[0][0][7][0]),
.cpatr_o_0_0_7_1_V(wire_cpatr_o[0][0][7][1]),
.cpatr_o_0_0_8_0_V(wire_cpatr_o[0][0][8][0]),
.cpatr_o_0_0_8_1_V(wire_cpatr_o[0][0][8][1]),
.cpatr_o_0_1_0_0_V(wire_cpatr_o[0][1][0][0]),
.cpatr_o_0_1_0_1_V(wire_cpatr_o[0][1][0][1]),
.cpatr_o_0_1_1_0_V(wire_cpatr_o[0][1][1][0]),
.cpatr_o_0_1_1_1_V(wire_cpatr_o[0][1][1][1]),
.cpatr_o_0_1_2_0_V(wire_cpatr_o[0][1][2][0]),
.cpatr_o_0_1_2_1_V(wire_cpatr_o[0][1][2][1]),
.cpatr_o_0_1_3_0_V(wire_cpatr_o[0][1][3][0]),
.cpatr_o_0_1_3_1_V(wire_cpatr_o[0][1][3][1]),
.cpatr_o_0_1_4_0_V(wire_cpatr_o[0][1][4][0]),
.cpatr_o_0_1_4_1_V(wire_cpatr_o[0][1][4][1]),
.cpatr_o_0_1_5_0_V(wire_cpatr_o[0][1][5][0]),
.cpatr_o_0_1_5_1_V(wire_cpatr_o[0][1][5][1]),
.cpatr_o_0_1_6_0_V(wire_cpatr_o[0][1][6][0]),
.cpatr_o_0_1_6_1_V(wire_cpatr_o[0][1][6][1]),
.cpatr_o_0_1_7_0_V(wire_cpatr_o[0][1][7][0]),
.cpatr_o_0_1_7_1_V(wire_cpatr_o[0][1][7][1]),
.cpatr_o_0_1_8_0_V(wire_cpatr_o[0][1][8][0]),
.cpatr_o_0_1_8_1_V(wire_cpatr_o[0][1][8][1]),
.cpatr_o_0_2_0_0_V(wire_cpatr_o[0][2][0][0]),
.cpatr_o_0_2_0_1_V(wire_cpatr_o[0][2][0][1]),
.cpatr_o_0_2_1_0_V(wire_cpatr_o[0][2][1][0]),
.cpatr_o_0_2_1_1_V(wire_cpatr_o[0][2][1][1]),
.cpatr_o_0_2_2_0_V(wire_cpatr_o[0][2][2][0]),
.cpatr_o_0_2_2_1_V(wire_cpatr_o[0][2][2][1]),
.cpatr_o_0_2_3_0_V(wire_cpatr_o[0][2][3][0]),
.cpatr_o_0_2_3_1_V(wire_cpatr_o[0][2][3][1]),
.cpatr_o_0_2_4_0_V(wire_cpatr_o[0][2][4][0]),
.cpatr_o_0_2_4_1_V(wire_cpatr_o[0][2][4][1]),
.cpatr_o_0_2_5_0_V(wire_cpatr_o[0][2][5][0]),
.cpatr_o_0_2_5_1_V(wire_cpatr_o[0][2][5][1]),
.cpatr_o_0_2_6_0_V(wire_cpatr_o[0][2][6][0]),
.cpatr_o_0_2_6_1_V(wire_cpatr_o[0][2][6][1]),
.cpatr_o_0_2_7_0_V(wire_cpatr_o[0][2][7][0]),
.cpatr_o_0_2_7_1_V(wire_cpatr_o[0][2][7][1]),
.cpatr_o_0_2_8_0_V(wire_cpatr_o[0][2][8][0]),
.cpatr_o_0_2_8_1_V(wire_cpatr_o[0][2][8][1]),
.cpatr_o_0_3_0_0_V(wire_cpatr_o[0][3][0][0]),
.cpatr_o_0_3_0_1_V(wire_cpatr_o[0][3][0][1]),
.cpatr_o_0_3_1_0_V(wire_cpatr_o[0][3][1][0]),
.cpatr_o_0_3_1_1_V(wire_cpatr_o[0][3][1][1]),
.cpatr_o_0_3_2_0_V(wire_cpatr_o[0][3][2][0]),
.cpatr_o_0_3_2_1_V(wire_cpatr_o[0][3][2][1]),
.cpatr_o_0_3_3_0_V(wire_cpatr_o[0][3][3][0]),
.cpatr_o_0_3_3_1_V(wire_cpatr_o[0][3][3][1]),
.cpatr_o_0_3_4_0_V(wire_cpatr_o[0][3][4][0]),
.cpatr_o_0_3_4_1_V(wire_cpatr_o[0][3][4][1]),
.cpatr_o_0_3_5_0_V(wire_cpatr_o[0][3][5][0]),
.cpatr_o_0_3_5_1_V(wire_cpatr_o[0][3][5][1]),
.cpatr_o_0_3_6_0_V(wire_cpatr_o[0][3][6][0]),
.cpatr_o_0_3_6_1_V(wire_cpatr_o[0][3][6][1]),
.cpatr_o_0_3_7_0_V(wire_cpatr_o[0][3][7][0]),
.cpatr_o_0_3_7_1_V(wire_cpatr_o[0][3][7][1]),
.cpatr_o_0_3_8_0_V(wire_cpatr_o[0][3][8][0]),
.cpatr_o_0_3_8_1_V(wire_cpatr_o[0][3][8][1]),
.cpatr_o_0_4_0_0_V(wire_cpatr_o[0][4][0][0]),
.cpatr_o_0_4_0_1_V(wire_cpatr_o[0][4][0][1]),
.cpatr_o_0_4_1_0_V(wire_cpatr_o[0][4][1][0]),
.cpatr_o_0_4_1_1_V(wire_cpatr_o[0][4][1][1]),
.cpatr_o_0_4_2_0_V(wire_cpatr_o[0][4][2][0]),
.cpatr_o_0_4_2_1_V(wire_cpatr_o[0][4][2][1]),
.cpatr_o_0_4_3_0_V(wire_cpatr_o[0][4][3][0]),
.cpatr_o_0_4_3_1_V(wire_cpatr_o[0][4][3][1]),
.cpatr_o_0_4_4_0_V(wire_cpatr_o[0][4][4][0]),
.cpatr_o_0_4_4_1_V(wire_cpatr_o[0][4][4][1]),
.cpatr_o_0_4_5_0_V(wire_cpatr_o[0][4][5][0]),
.cpatr_o_0_4_5_1_V(wire_cpatr_o[0][4][5][1]),
.cpatr_o_0_4_6_0_V(wire_cpatr_o[0][4][6][0]),
.cpatr_o_0_4_6_1_V(wire_cpatr_o[0][4][6][1]),
.cpatr_o_0_4_7_0_V(wire_cpatr_o[0][4][7][0]),
.cpatr_o_0_4_7_1_V(wire_cpatr_o[0][4][7][1]),
.cpatr_o_0_4_8_0_V(wire_cpatr_o[0][4][8][0]),
.cpatr_o_0_4_8_1_V(wire_cpatr_o[0][4][8][1]),
.cpatr_o_0_5_0_0_V(wire_cpatr_o[0][5][0][0]),
.cpatr_o_0_5_0_1_V(wire_cpatr_o[0][5][0][1]),
.cpatr_o_0_5_1_0_V(wire_cpatr_o[0][5][1][0]),
.cpatr_o_0_5_1_1_V(wire_cpatr_o[0][5][1][1]),
.cpatr_o_0_5_2_0_V(wire_cpatr_o[0][5][2][0]),
.cpatr_o_0_5_2_1_V(wire_cpatr_o[0][5][2][1]),
.cpatr_o_0_5_3_0_V(wire_cpatr_o[0][5][3][0]),
.cpatr_o_0_5_3_1_V(wire_cpatr_o[0][5][3][1]),
.cpatr_o_0_5_4_0_V(wire_cpatr_o[0][5][4][0]),
.cpatr_o_0_5_4_1_V(wire_cpatr_o[0][5][4][1]),
.cpatr_o_0_5_5_0_V(wire_cpatr_o[0][5][5][0]),
.cpatr_o_0_5_5_1_V(wire_cpatr_o[0][5][5][1]),
.cpatr_o_0_5_6_0_V(wire_cpatr_o[0][5][6][0]),
.cpatr_o_0_5_6_1_V(wire_cpatr_o[0][5][6][1]),
.cpatr_o_0_5_7_0_V(wire_cpatr_o[0][5][7][0]),
.cpatr_o_0_5_7_1_V(wire_cpatr_o[0][5][7][1]),
.cpatr_o_0_5_8_0_V(wire_cpatr_o[0][5][8][0]),
.cpatr_o_0_5_8_1_V(wire_cpatr_o[0][5][8][1]),
.ph_o_0_0_0_0_V(wire_ph_o[0][0][0][0]),
.ph_o_0_0_0_1_V(wire_ph_o[0][0][0][1]),
.ph_o_0_0_1_0_V(wire_ph_o[0][0][1][0]),
.ph_o_0_0_1_1_V(wire_ph_o[0][0][1][1]),
.ph_o_0_0_2_0_V(wire_ph_o[0][0][2][0]),
.ph_o_0_0_2_1_V(wire_ph_o[0][0][2][1]),
.ph_o_0_0_3_0_V(wire_ph_o[0][0][3][0]),
.ph_o_0_0_3_1_V(wire_ph_o[0][0][3][1]),
.ph_o_0_0_4_0_V(wire_ph_o[0][0][4][0]),
.ph_o_0_0_4_1_V(wire_ph_o[0][0][4][1]),
.ph_o_0_0_5_0_V(wire_ph_o[0][0][5][0]),
.ph_o_0_0_5_1_V(wire_ph_o[0][0][5][1]),
.ph_o_0_0_6_0_V(wire_ph_o[0][0][6][0]),
.ph_o_0_0_6_1_V(wire_ph_o[0][0][6][1]),
.ph_o_0_0_7_0_V(wire_ph_o[0][0][7][0]),
.ph_o_0_0_7_1_V(wire_ph_o[0][0][7][1]),
.ph_o_0_0_8_0_V(wire_ph_o[0][0][8][0]),
.ph_o_0_0_8_1_V(wire_ph_o[0][0][8][1]),
.ph_o_0_1_0_0_V(wire_ph_o[0][1][0][0]),
.ph_o_0_1_0_1_V(wire_ph_o[0][1][0][1]),
.ph_o_0_1_1_0_V(wire_ph_o[0][1][1][0]),
.ph_o_0_1_1_1_V(wire_ph_o[0][1][1][1]),
.ph_o_0_1_2_0_V(wire_ph_o[0][1][2][0]),
.ph_o_0_1_2_1_V(wire_ph_o[0][1][2][1]),
.ph_o_0_1_3_0_V(wire_ph_o[0][1][3][0]),
.ph_o_0_1_3_1_V(wire_ph_o[0][1][3][1]),
.ph_o_0_1_4_0_V(wire_ph_o[0][1][4][0]),
.ph_o_0_1_4_1_V(wire_ph_o[0][1][4][1]),
.ph_o_0_1_5_0_V(wire_ph_o[0][1][5][0]),
.ph_o_0_1_5_1_V(wire_ph_o[0][1][5][1]),
.ph_o_0_1_6_0_V(wire_ph_o[0][1][6][0]),
.ph_o_0_1_6_1_V(wire_ph_o[0][1][6][1]),
.ph_o_0_1_7_0_V(wire_ph_o[0][1][7][0]),
.ph_o_0_1_7_1_V(wire_ph_o[0][1][7][1]),
.ph_o_0_1_8_0_V(wire_ph_o[0][1][8][0]),
.ph_o_0_1_8_1_V(wire_ph_o[0][1][8][1]),
.ph_o_0_2_0_0_V(wire_ph_o[0][2][0][0]),
.ph_o_0_2_0_1_V(wire_ph_o[0][2][0][1]),
.ph_o_0_2_1_0_V(wire_ph_o[0][2][1][0]),
.ph_o_0_2_1_1_V(wire_ph_o[0][2][1][1]),
.ph_o_0_2_2_0_V(wire_ph_o[0][2][2][0]),
.ph_o_0_2_2_1_V(wire_ph_o[0][2][2][1]),
.ph_o_0_2_3_0_V(wire_ph_o[0][2][3][0]),
.ph_o_0_2_3_1_V(wire_ph_o[0][2][3][1]),
.ph_o_0_2_4_0_V(wire_ph_o[0][2][4][0]),
.ph_o_0_2_4_1_V(wire_ph_o[0][2][4][1]),
.ph_o_0_2_5_0_V(wire_ph_o[0][2][5][0]),
.ph_o_0_2_5_1_V(wire_ph_o[0][2][5][1]),
.ph_o_0_2_6_0_V(wire_ph_o[0][2][6][0]),
.ph_o_0_2_6_1_V(wire_ph_o[0][2][6][1]),
.ph_o_0_2_7_0_V(wire_ph_o[0][2][7][0]),
.ph_o_0_2_7_1_V(wire_ph_o[0][2][7][1]),
.ph_o_0_2_8_0_V(wire_ph_o[0][2][8][0]),
.ph_o_0_2_8_1_V(wire_ph_o[0][2][8][1]),
.ph_o_0_3_0_0_V(wire_ph_o[0][3][0][0]),
.ph_o_0_3_0_1_V(wire_ph_o[0][3][0][1]),
.ph_o_0_3_1_0_V(wire_ph_o[0][3][1][0]),
.ph_o_0_3_1_1_V(wire_ph_o[0][3][1][1]),
.ph_o_0_3_2_0_V(wire_ph_o[0][3][2][0]),
.ph_o_0_3_2_1_V(wire_ph_o[0][3][2][1]),
.ph_o_0_3_3_0_V(wire_ph_o[0][3][3][0]),
.ph_o_0_3_3_1_V(wire_ph_o[0][3][3][1]),
.ph_o_0_3_4_0_V(wire_ph_o[0][3][4][0]),
.ph_o_0_3_4_1_V(wire_ph_o[0][3][4][1]),
.ph_o_0_3_5_0_V(wire_ph_o[0][3][5][0]),
.ph_o_0_3_5_1_V(wire_ph_o[0][3][5][1]),
.ph_o_0_3_6_0_V(wire_ph_o[0][3][6][0]),
.ph_o_0_3_6_1_V(wire_ph_o[0][3][6][1]),
.ph_o_0_3_7_0_V(wire_ph_o[0][3][7][0]),
.ph_o_0_3_7_1_V(wire_ph_o[0][3][7][1]),
.ph_o_0_3_8_0_V(wire_ph_o[0][3][8][0]),
.ph_o_0_3_8_1_V(wire_ph_o[0][3][8][1]),
.ph_o_0_4_0_0_V(wire_ph_o[0][4][0][0]),
.ph_o_0_4_0_1_V(wire_ph_o[0][4][0][1]),
.ph_o_0_4_1_0_V(wire_ph_o[0][4][1][0]),
.ph_o_0_4_1_1_V(wire_ph_o[0][4][1][1]),
.ph_o_0_4_2_0_V(wire_ph_o[0][4][2][0]),
.ph_o_0_4_2_1_V(wire_ph_o[0][4][2][1]),
.ph_o_0_4_3_0_V(wire_ph_o[0][4][3][0]),
.ph_o_0_4_3_1_V(wire_ph_o[0][4][3][1]),
.ph_o_0_4_4_0_V(wire_ph_o[0][4][4][0]),
.ph_o_0_4_4_1_V(wire_ph_o[0][4][4][1]),
.ph_o_0_4_5_0_V(wire_ph_o[0][4][5][0]),
.ph_o_0_4_5_1_V(wire_ph_o[0][4][5][1]),
.ph_o_0_4_6_0_V(wire_ph_o[0][4][6][0]),
.ph_o_0_4_6_1_V(wire_ph_o[0][4][6][1]),
.ph_o_0_4_7_0_V(wire_ph_o[0][4][7][0]),
.ph_o_0_4_7_1_V(wire_ph_o[0][4][7][1]),
.ph_o_0_4_8_0_V(wire_ph_o[0][4][8][0]),
.ph_o_0_4_8_1_V(wire_ph_o[0][4][8][1]),
.ph_o_0_5_0_0_V(wire_ph_o[0][5][0][0]),
.ph_o_0_5_0_1_V(wire_ph_o[0][5][0][1]),
.ph_o_0_5_1_0_V(wire_ph_o[0][5][1][0]),
.ph_o_0_5_1_1_V(wire_ph_o[0][5][1][1]),
.ph_o_0_5_2_0_V(wire_ph_o[0][5][2][0]),
.ph_o_0_5_2_1_V(wire_ph_o[0][5][2][1]),
.ph_o_0_5_3_0_V(wire_ph_o[0][5][3][0]),
.ph_o_0_5_3_1_V(wire_ph_o[0][5][3][1]),
.ph_o_0_5_4_0_V(wire_ph_o[0][5][4][0]),
.ph_o_0_5_4_1_V(wire_ph_o[0][5][4][1]),
.ph_o_0_5_5_0_V(wire_ph_o[0][5][5][0]),
.ph_o_0_5_5_1_V(wire_ph_o[0][5][5][1]),
.ph_o_0_5_6_0_V(wire_ph_o[0][5][6][0]),
.ph_o_0_5_6_1_V(wire_ph_o[0][5][6][1]),
.ph_o_0_5_7_0_V(wire_ph_o[0][5][7][0]),
.ph_o_0_5_7_1_V(wire_ph_o[0][5][7][1]),
.ph_o_0_5_8_0_V(wire_ph_o[0][5][8][0]),
.ph_o_0_5_8_1_V(wire_ph_o[0][5][8][1]),
.th11_o_0_0_0_0_V(wire_th11_o[0][0][0][0]),
.th11_o_0_0_0_1_V(wire_th11_o[0][0][0][1]),
.th11_o_0_0_1_0_V(wire_th11_o[0][0][1][0]),
.th11_o_0_0_1_1_V(wire_th11_o[0][0][1][1]),
.th11_o_0_0_2_0_V(wire_th11_o[0][0][2][0]),
.th11_o_0_0_2_1_V(wire_th11_o[0][0][2][1]),
.th11_o_0_0_3_0_V(wire_th11_o[0][0][3][0]),
.th11_o_0_0_3_1_V(wire_th11_o[0][0][3][1]),
.th11_o_0_0_4_0_V(wire_th11_o[0][0][4][0]),
.th11_o_0_0_4_1_V(wire_th11_o[0][0][4][1]),
.th11_o_0_0_5_0_V(wire_th11_o[0][0][5][0]),
.th11_o_0_0_5_1_V(wire_th11_o[0][0][5][1]),
.th11_o_0_0_6_0_V(wire_th11_o[0][0][6][0]),
.th11_o_0_0_6_1_V(wire_th11_o[0][0][6][1]),
.th11_o_0_0_7_0_V(wire_th11_o[0][0][7][0]),
.th11_o_0_0_7_1_V(wire_th11_o[0][0][7][1]),
.th11_o_0_0_8_0_V(wire_th11_o[0][0][8][0]),
.th11_o_0_0_8_1_V(wire_th11_o[0][0][8][1]),
.th11_o_0_1_0_0_V(wire_th11_o[0][1][0][0]),
.th11_o_0_1_0_1_V(wire_th11_o[0][1][0][1]),
.th11_o_0_1_1_0_V(wire_th11_o[0][1][1][0]),
.th11_o_0_1_1_1_V(wire_th11_o[0][1][1][1]),
.th11_o_0_1_2_0_V(wire_th11_o[0][1][2][0]),
.th11_o_0_1_2_1_V(wire_th11_o[0][1][2][1]),
.th11_o_0_1_3_0_V(wire_th11_o[0][1][3][0]),
.th11_o_0_1_3_1_V(wire_th11_o[0][1][3][1]),
.th11_o_0_1_4_0_V(wire_th11_o[0][1][4][0]),
.th11_o_0_1_4_1_V(wire_th11_o[0][1][4][1]),
.th11_o_0_1_5_0_V(wire_th11_o[0][1][5][0]),
.th11_o_0_1_5_1_V(wire_th11_o[0][1][5][1]),
.th11_o_0_1_6_0_V(wire_th11_o[0][1][6][0]),
.th11_o_0_1_6_1_V(wire_th11_o[0][1][6][1]),
.th11_o_0_1_7_0_V(wire_th11_o[0][1][7][0]),
.th11_o_0_1_7_1_V(wire_th11_o[0][1][7][1]),
.th11_o_0_1_8_0_V(wire_th11_o[0][1][8][0]),
.th11_o_0_1_8_1_V(wire_th11_o[0][1][8][1]),
.th11_o_0_2_0_0_V(wire_th11_o[0][2][0][0]),
.th11_o_0_2_0_1_V(wire_th11_o[0][2][0][1]),
.th11_o_0_2_1_0_V(wire_th11_o[0][2][1][0]),
.th11_o_0_2_1_1_V(wire_th11_o[0][2][1][1]),
.th11_o_0_2_2_0_V(wire_th11_o[0][2][2][0]),
.th11_o_0_2_2_1_V(wire_th11_o[0][2][2][1]),
.th11_o_0_2_3_0_V(wire_th11_o[0][2][3][0]),
.th11_o_0_2_3_1_V(wire_th11_o[0][2][3][1]),
.th11_o_0_2_4_0_V(wire_th11_o[0][2][4][0]),
.th11_o_0_2_4_1_V(wire_th11_o[0][2][4][1]),
.th11_o_0_2_5_0_V(wire_th11_o[0][2][5][0]),
.th11_o_0_2_5_1_V(wire_th11_o[0][2][5][1]),
.th11_o_0_2_6_0_V(wire_th11_o[0][2][6][0]),
.th11_o_0_2_6_1_V(wire_th11_o[0][2][6][1]),
.th11_o_0_2_7_0_V(wire_th11_o[0][2][7][0]),
.th11_o_0_2_7_1_V(wire_th11_o[0][2][7][1]),
.th11_o_0_2_8_0_V(wire_th11_o[0][2][8][0]),
.th11_o_0_2_8_1_V(wire_th11_o[0][2][8][1]),
.th11_o_0_3_0_0_V(wire_th11_o[0][3][0][0]),
.th11_o_0_3_0_1_V(wire_th11_o[0][3][0][1]),
.th11_o_0_3_1_0_V(wire_th11_o[0][3][1][0]),
.th11_o_0_3_1_1_V(wire_th11_o[0][3][1][1]),
.th11_o_0_3_2_0_V(wire_th11_o[0][3][2][0]),
.th11_o_0_3_2_1_V(wire_th11_o[0][3][2][1]),
.th11_o_0_3_3_0_V(wire_th11_o[0][3][3][0]),
.th11_o_0_3_3_1_V(wire_th11_o[0][3][3][1]),
.th11_o_0_3_4_0_V(wire_th11_o[0][3][4][0]),
.th11_o_0_3_4_1_V(wire_th11_o[0][3][4][1]),
.th11_o_0_3_5_0_V(wire_th11_o[0][3][5][0]),
.th11_o_0_3_5_1_V(wire_th11_o[0][3][5][1]),
.th11_o_0_3_6_0_V(wire_th11_o[0][3][6][0]),
.th11_o_0_3_6_1_V(wire_th11_o[0][3][6][1]),
.th11_o_0_3_7_0_V(wire_th11_o[0][3][7][0]),
.th11_o_0_3_7_1_V(wire_th11_o[0][3][7][1]),
.th11_o_0_3_8_0_V(wire_th11_o[0][3][8][0]),
.th11_o_0_3_8_1_V(wire_th11_o[0][3][8][1]),
.th11_o_0_4_0_0_V(wire_th11_o[0][4][0][0]),
.th11_o_0_4_0_1_V(wire_th11_o[0][4][0][1]),
.th11_o_0_4_1_0_V(wire_th11_o[0][4][1][0]),
.th11_o_0_4_1_1_V(wire_th11_o[0][4][1][1]),
.th11_o_0_4_2_0_V(wire_th11_o[0][4][2][0]),
.th11_o_0_4_2_1_V(wire_th11_o[0][4][2][1]),
.th11_o_0_4_3_0_V(wire_th11_o[0][4][3][0]),
.th11_o_0_4_3_1_V(wire_th11_o[0][4][3][1]),
.th11_o_0_4_4_0_V(wire_th11_o[0][4][4][0]),
.th11_o_0_4_4_1_V(wire_th11_o[0][4][4][1]),
.th11_o_0_4_5_0_V(wire_th11_o[0][4][5][0]),
.th11_o_0_4_5_1_V(wire_th11_o[0][4][5][1]),
.th11_o_0_4_6_0_V(wire_th11_o[0][4][6][0]),
.th11_o_0_4_6_1_V(wire_th11_o[0][4][6][1]),
.th11_o_0_4_7_0_V(wire_th11_o[0][4][7][0]),
.th11_o_0_4_7_1_V(wire_th11_o[0][4][7][1]),
.th11_o_0_4_8_0_V(wire_th11_o[0][4][8][0]),
.th11_o_0_4_8_1_V(wire_th11_o[0][4][8][1]),
.th11_o_0_5_0_0_V(wire_th11_o[0][5][0][0]),
.th11_o_0_5_0_1_V(wire_th11_o[0][5][0][1]),
.th11_o_0_5_1_0_V(wire_th11_o[0][5][1][0]),
.th11_o_0_5_1_1_V(wire_th11_o[0][5][1][1]),
.th11_o_0_5_2_0_V(wire_th11_o[0][5][2][0]),
.th11_o_0_5_2_1_V(wire_th11_o[0][5][2][1]),
.th11_o_0_5_3_0_V(wire_th11_o[0][5][3][0]),
.th11_o_0_5_3_1_V(wire_th11_o[0][5][3][1]),
.th11_o_0_5_4_0_V(wire_th11_o[0][5][4][0]),
.th11_o_0_5_4_1_V(wire_th11_o[0][5][4][1]),
.th11_o_0_5_5_0_V(wire_th11_o[0][5][5][0]),
.th11_o_0_5_5_1_V(wire_th11_o[0][5][5][1]),
.th11_o_0_5_6_0_V(wire_th11_o[0][5][6][0]),
.th11_o_0_5_6_1_V(wire_th11_o[0][5][6][1]),
.th11_o_0_5_7_0_V(wire_th11_o[0][5][7][0]),
.th11_o_0_5_7_1_V(wire_th11_o[0][5][7][1]),
.th11_o_0_5_8_0_V(wire_th11_o[0][5][8][0]),
.th11_o_0_5_8_1_V(wire_th11_o[0][5][8][1]),
.th_o_0_0_0_0_V(wire_th_o[0][0][0][0]),
.th_o_0_0_0_1_V(wire_th_o[0][0][0][1]),
.th_o_0_0_0_2_V(wire_th_o[0][0][0][2]),
.th_o_0_0_0_3_V(wire_th_o[0][0][0][3]),
.th_o_0_0_1_0_V(wire_th_o[0][0][1][0]),
.th_o_0_0_1_1_V(wire_th_o[0][0][1][1]),
.th_o_0_0_1_2_V(wire_th_o[0][0][1][2]),
.th_o_0_0_1_3_V(wire_th_o[0][0][1][3]),
.th_o_0_0_2_0_V(wire_th_o[0][0][2][0]),
.th_o_0_0_2_1_V(wire_th_o[0][0][2][1]),
.th_o_0_0_2_2_V(wire_th_o[0][0][2][2]),
.th_o_0_0_2_3_V(wire_th_o[0][0][2][3]),
.th_o_0_1_0_0_V(wire_th_o[0][1][0][0]),
.th_o_0_1_0_1_V(wire_th_o[0][1][0][1]),
.th_o_0_1_0_2_V(wire_th_o[0][1][0][2]),
.th_o_0_1_0_3_V(wire_th_o[0][1][0][3]),
.th_o_0_1_1_0_V(wire_th_o[0][1][1][0]),
.th_o_0_1_1_1_V(wire_th_o[0][1][1][1]),
.th_o_0_1_1_2_V(wire_th_o[0][1][1][2]),
.th_o_0_1_1_3_V(wire_th_o[0][1][1][3]),
.th_o_0_1_2_0_V(wire_th_o[0][1][2][0]),
.th_o_0_1_2_1_V(wire_th_o[0][1][2][1]),
.th_o_0_1_2_2_V(wire_th_o[0][1][2][2]),
.th_o_0_1_2_3_V(wire_th_o[0][1][2][3]),
.th_o_0_2_0_0_V(wire_th_o[0][2][0][0]),
.th_o_0_2_0_1_V(wire_th_o[0][2][0][1]),
.th_o_0_2_0_2_V(wire_th_o[0][2][0][2]),
.th_o_0_2_0_3_V(wire_th_o[0][2][0][3]),
.th_o_0_2_1_0_V(wire_th_o[0][2][1][0]),
.th_o_0_2_1_1_V(wire_th_o[0][2][1][1]),
.th_o_0_2_1_2_V(wire_th_o[0][2][1][2]),
.th_o_0_2_1_3_V(wire_th_o[0][2][1][3]),
.th_o_0_2_2_0_V(wire_th_o[0][2][2][0]),
.th_o_0_2_2_1_V(wire_th_o[0][2][2][1]),
.th_o_0_2_2_2_V(wire_th_o[0][2][2][2]),
.th_o_0_2_2_3_V(wire_th_o[0][2][2][3]),
.phzvl_o_0_0_0_V(wire_phzvl_o[0][0][0]),
.phzvl_o_0_0_1_V(wire_phzvl_o[0][0][1]),
.phzvl_o_0_0_2_V(wire_phzvl_o[0][0][2]),
.phzvl_o_0_0_3_V(wire_phzvl_o[0][0][3]),
.phzvl_o_0_0_4_V(wire_phzvl_o[0][0][4]),
.phzvl_o_0_0_5_V(wire_phzvl_o[0][0][5]),
.phzvl_o_0_0_6_V(wire_phzvl_o[0][0][6]),
.phzvl_o_0_0_7_V(wire_phzvl_o[0][0][7]),
.phzvl_o_0_0_8_V(wire_phzvl_o[0][0][8]),
.phzvl_o_0_1_0_V(wire_phzvl_o[0][1][0]),
.phzvl_o_0_1_1_V(wire_phzvl_o[0][1][1]),
.phzvl_o_0_1_2_V(wire_phzvl_o[0][1][2]),
.phzvl_o_0_1_3_V(wire_phzvl_o[0][1][3]),
.phzvl_o_0_1_4_V(wire_phzvl_o[0][1][4]),
.phzvl_o_0_1_5_V(wire_phzvl_o[0][1][5]),
.phzvl_o_0_1_6_V(wire_phzvl_o[0][1][6]),
.phzvl_o_0_1_7_V(wire_phzvl_o[0][1][7]),
.phzvl_o_0_1_8_V(wire_phzvl_o[0][1][8]),
.phzvl_o_0_2_0_V(wire_phzvl_o[0][2][0]),
.phzvl_o_0_2_1_V(wire_phzvl_o[0][2][1]),
.phzvl_o_0_2_2_V(wire_phzvl_o[0][2][2]),
.phzvl_o_0_2_3_V(wire_phzvl_o[0][2][3]),
.phzvl_o_0_2_4_V(wire_phzvl_o[0][2][4]),
.phzvl_o_0_2_5_V(wire_phzvl_o[0][2][5]),
.phzvl_o_0_2_6_V(wire_phzvl_o[0][2][6]),
.phzvl_o_0_2_7_V(wire_phzvl_o[0][2][7]),
.phzvl_o_0_2_8_V(wire_phzvl_o[0][2][8]),
.phzvl_o_0_3_0_V(wire_phzvl_o[0][3][0]),
.phzvl_o_0_3_1_V(wire_phzvl_o[0][3][1]),
.phzvl_o_0_3_2_V(wire_phzvl_o[0][3][2]),
.phzvl_o_0_3_3_V(wire_phzvl_o[0][3][3]),
.phzvl_o_0_3_4_V(wire_phzvl_o[0][3][4]),
.phzvl_o_0_3_5_V(wire_phzvl_o[0][3][5]),
.phzvl_o_0_3_6_V(wire_phzvl_o[0][3][6]),
.phzvl_o_0_3_7_V(wire_phzvl_o[0][3][7]),
.phzvl_o_0_3_8_V(wire_phzvl_o[0][3][8]),
.phzvl_o_0_4_0_V(wire_phzvl_o[0][4][0]),
.phzvl_o_0_4_1_V(wire_phzvl_o[0][4][1]),
.phzvl_o_0_4_2_V(wire_phzvl_o[0][4][2]),
.phzvl_o_0_4_3_V(wire_phzvl_o[0][4][3]),
.phzvl_o_0_4_4_V(wire_phzvl_o[0][4][4]),
.phzvl_o_0_4_5_V(wire_phzvl_o[0][4][5]),
.phzvl_o_0_4_6_V(wire_phzvl_o[0][4][6]),
.phzvl_o_0_4_7_V(wire_phzvl_o[0][4][7]),
.phzvl_o_0_4_8_V(wire_phzvl_o[0][4][8]),
.phzvl_o_0_5_0_V(wire_phzvl_o[0][5][0]),
.phzvl_o_0_5_1_V(wire_phzvl_o[0][5][1]),
.phzvl_o_0_5_2_V(wire_phzvl_o[0][5][2]),
.phzvl_o_0_5_3_V(wire_phzvl_o[0][5][3]),
.phzvl_o_0_5_4_V(wire_phzvl_o[0][5][4]),
.phzvl_o_0_5_5_V(wire_phzvl_o[0][5][5]),
.phzvl_o_0_5_6_V(wire_phzvl_o[0][5][6]),
.phzvl_o_0_5_7_V(wire_phzvl_o[0][5][7]),
.phzvl_o_0_5_8_V(wire_phzvl_o[0][5][8]),
.phzvl_o_0_6_0_V(wire_phzvl_o[0][6][0]),
.phzvl_o_0_6_1_V(wire_phzvl_o[0][6][1]),
.phzvl_o_0_6_2_V(wire_phzvl_o[0][6][2]),
.phzvl_o_0_6_3_V(wire_phzvl_o[0][6][3]),
.phzvl_o_0_6_4_V(wire_phzvl_o[0][6][4]),
.phzvl_o_0_6_5_V(wire_phzvl_o[0][6][5]),
.phzvl_o_0_6_6_V(wire_phzvl_o[0][6][6]),
.phzvl_o_0_6_7_V(wire_phzvl_o[0][6][7]),
.phzvl_o_0_6_8_V(wire_phzvl_o[0][6][8]),
.phzvl_o_0_7_0_V(wire_phzvl_o[0][7][0]),
.phzvl_o_0_7_1_V(wire_phzvl_o[0][7][1]),
.phzvl_o_0_7_2_V(wire_phzvl_o[0][7][2]),
.phzvl_o_0_7_3_V(wire_phzvl_o[0][7][3]),
.phzvl_o_0_7_4_V(wire_phzvl_o[0][7][4]),
.phzvl_o_0_7_5_V(wire_phzvl_o[0][7][5]),
.phzvl_o_0_7_6_V(wire_phzvl_o[0][7][6]),
.phzvl_o_0_7_7_V(wire_phzvl_o[0][7][7]),
.phzvl_o_0_7_8_V(wire_phzvl_o[0][7][8]),
.phzvl_o_0_8_0_V(wire_phzvl_o[0][8][0]),
.phzvl_o_0_8_1_V(wire_phzvl_o[0][8][1]),
.phzvl_o_0_8_2_V(wire_phzvl_o[0][8][2]),
.phzvl_o_0_8_3_V(wire_phzvl_o[0][8][3]),
.phzvl_o_0_8_4_V(wire_phzvl_o[0][8][4]),
.phzvl_o_0_8_5_V(wire_phzvl_o[0][8][5]),
.phzvl_o_0_8_6_V(wire_phzvl_o[0][8][6]),
.phzvl_o_0_8_7_V(wire_phzvl_o[0][8][7]),
.phzvl_o_0_8_8_V(wire_phzvl_o[0][8][8]),
.phzvl_o_0_9_0_V(wire_phzvl_o[0][9][0]),
.phzvl_o_0_9_1_V(wire_phzvl_o[0][9][1]),
.phzvl_o_0_9_2_V(wire_phzvl_o[0][9][2]),
.phzvl_o_0_9_3_V(wire_phzvl_o[0][9][3]),
.phzvl_o_0_9_4_V(wire_phzvl_o[0][9][4]),
.phzvl_o_0_9_5_V(wire_phzvl_o[0][9][5]),
.phzvl_o_0_9_6_V(wire_phzvl_o[0][9][6]),
.phzvl_o_0_9_7_V(wire_phzvl_o[0][9][7]),
.phzvl_o_0_9_8_V(wire_phzvl_o[0][9][8]),
.phzvl_o_0_10_0_V(wire_phzvl_o[0][10][0]),
.phzvl_o_0_10_1_V(wire_phzvl_o[0][10][1]),
.phzvl_o_0_10_2_V(wire_phzvl_o[0][10][2]),
.phzvl_o_0_10_3_V(wire_phzvl_o[0][10][3]),
.phzvl_o_0_10_4_V(wire_phzvl_o[0][10][4]),
.phzvl_o_0_10_5_V(wire_phzvl_o[0][10][5]),
.phzvl_o_0_10_6_V(wire_phzvl_o[0][10][6]),
.phzvl_o_0_10_7_V(wire_phzvl_o[0][10][7]),
.phzvl_o_0_10_8_V(wire_phzvl_o[0][10][8]),
.phzvl_o_0_11_0_V(wire_phzvl_o[0][11][0]),
.phzvl_o_0_11_1_V(wire_phzvl_o[0][11][1]),
.phzvl_o_0_11_2_V(wire_phzvl_o[0][11][2]),
.phzvl_o_0_11_3_V(wire_phzvl_o[0][11][3]),
.phzvl_o_0_11_4_V(wire_phzvl_o[0][11][4]),
.phzvl_o_0_11_5_V(wire_phzvl_o[0][11][5]),
.phzvl_o_0_11_6_V(wire_phzvl_o[0][11][6]),
.phzvl_o_0_11_7_V(wire_phzvl_o[0][11][7]),
.phzvl_o_0_11_8_V(wire_phzvl_o[0][11][8]),
.phzvl_o_0_12_0_V(wire_phzvl_o[0][12][0]),
.phzvl_o_0_12_1_V(wire_phzvl_o[0][12][1]),
.phzvl_o_0_12_2_V(wire_phzvl_o[0][12][2]),
.phzvl_o_0_12_3_V(wire_phzvl_o[0][12][3]),
.phzvl_o_0_12_4_V(wire_phzvl_o[0][12][4]),
.phzvl_o_0_12_5_V(wire_phzvl_o[0][12][5]),
.phzvl_o_0_12_6_V(wire_phzvl_o[0][12][6]),
.phzvl_o_0_12_7_V(wire_phzvl_o[0][12][7]),
.phzvl_o_0_12_8_V(wire_phzvl_o[0][12][8]),
.ph_hit_o_0_0_0_V(wire_ph_hit_o[0][0][0]),
.ph_hit_o_0_0_1_V(wire_ph_hit_o[0][0][1]),
.ph_hit_o_0_0_2_V(wire_ph_hit_o[0][0][2]),
.ph_hit_o_0_0_3_V(wire_ph_hit_o[0][0][3]),
.ph_hit_o_0_0_4_V(wire_ph_hit_o[0][0][4]),
.ph_hit_o_0_0_5_V(wire_ph_hit_o[0][0][5]),
.ph_hit_o_0_0_6_V(wire_ph_hit_o[0][0][6]),
.ph_hit_o_0_0_7_V(wire_ph_hit_o[0][0][7]),
.ph_hit_o_0_0_8_V(wire_ph_hit_o[0][0][8]),
.ph_hit_o_0_1_0_V(wire_ph_hit_o[0][1][0]),
.ph_hit_o_0_1_1_V(wire_ph_hit_o[0][1][1]),
.ph_hit_o_0_1_2_V(wire_ph_hit_o[0][1][2]),
.ph_hit_o_0_1_3_V(wire_ph_hit_o[0][1][3]),
.ph_hit_o_0_1_4_V(wire_ph_hit_o[0][1][4]),
.ph_hit_o_0_1_5_V(wire_ph_hit_o[0][1][5]),
.ph_hit_o_0_1_6_V(wire_ph_hit_o[0][1][6]),
.ph_hit_o_0_1_7_V(wire_ph_hit_o[0][1][7]),
.ph_hit_o_0_1_8_V(wire_ph_hit_o[0][1][8]),
.ph_hit_o_0_2_0_V(wire_ph_hit_o[0][2][0]),
.ph_hit_o_0_2_1_V(wire_ph_hit_o[0][2][1]),
.ph_hit_o_0_2_2_V(wire_ph_hit_o[0][2][2]),
.ph_hit_o_0_2_3_V(wire_ph_hit_o[0][2][3]),
.ph_hit_o_0_2_4_V(wire_ph_hit_o[0][2][4]),
.ph_hit_o_0_2_5_V(wire_ph_hit_o[0][2][5]),
.ph_hit_o_0_2_6_V(wire_ph_hit_o[0][2][6]),
.ph_hit_o_0_2_7_V(wire_ph_hit_o[0][2][7]),
.ph_hit_o_0_2_8_V(wire_ph_hit_o[0][2][8]),
.ph_hit_o_0_3_0_V(wire_ph_hit_o[0][3][0]),
.ph_hit_o_0_3_1_V(wire_ph_hit_o[0][3][1]),
.ph_hit_o_0_3_2_V(wire_ph_hit_o[0][3][2]),
.ph_hit_o_0_3_3_V(wire_ph_hit_o[0][3][3]),
.ph_hit_o_0_3_4_V(wire_ph_hit_o[0][3][4]),
.ph_hit_o_0_3_5_V(wire_ph_hit_o[0][3][5]),
.ph_hit_o_0_3_6_V(wire_ph_hit_o[0][3][6]),
.ph_hit_o_0_3_7_V(wire_ph_hit_o[0][3][7]),
.ph_hit_o_0_3_8_V(wire_ph_hit_o[0][3][8]),
.ph_hit_o_0_4_0_V(wire_ph_hit_o[0][4][0]),
.ph_hit_o_0_4_1_V(wire_ph_hit_o[0][4][1]),
.ph_hit_o_0_4_2_V(wire_ph_hit_o[0][4][2]),
.ph_hit_o_0_4_3_V(wire_ph_hit_o[0][4][3]),
.ph_hit_o_0_4_4_V(wire_ph_hit_o[0][4][4]),
.ph_hit_o_0_4_5_V(wire_ph_hit_o[0][4][5]),
.ph_hit_o_0_4_6_V(wire_ph_hit_o[0][4][6]),
.ph_hit_o_0_4_7_V(wire_ph_hit_o[0][4][7]),
.ph_hit_o_0_4_8_V(wire_ph_hit_o[0][4][8]),
.ph_hit_o_0_5_0_V(wire_ph_hit_o[0][5][0]),
.ph_hit_o_0_5_1_V(wire_ph_hit_o[0][5][1]),
.ph_hit_o_0_5_2_V(wire_ph_hit_o[0][5][2]),
.ph_hit_o_0_5_3_V(wire_ph_hit_o[0][5][3]),
.ph_hit_o_0_5_4_V(wire_ph_hit_o[0][5][4]),
.ph_hit_o_0_5_5_V(wire_ph_hit_o[0][5][5]),
.ph_hit_o_0_5_6_V(wire_ph_hit_o[0][5][6]),
.ph_hit_o_0_5_7_V(wire_ph_hit_o[0][5][7]),
.ph_hit_o_0_5_8_V(wire_ph_hit_o[0][5][8]),
.ph_hit_o_0_6_0_V(wire_ph_hit_o[0][6][0]),
.ph_hit_o_0_6_1_V(wire_ph_hit_o[0][6][1]),
.ph_hit_o_0_6_2_V(wire_ph_hit_o[0][6][2]),
.ph_hit_o_0_6_3_V(wire_ph_hit_o[0][6][3]),
.ph_hit_o_0_6_4_V(wire_ph_hit_o[0][6][4]),
.ph_hit_o_0_6_5_V(wire_ph_hit_o[0][6][5]),
.ph_hit_o_0_6_6_V(wire_ph_hit_o[0][6][6]),
.ph_hit_o_0_6_7_V(wire_ph_hit_o[0][6][7]),
.ph_hit_o_0_6_8_V(wire_ph_hit_o[0][6][8]),
.ph_hit_o_0_7_0_V(wire_ph_hit_o[0][7][0]),
.ph_hit_o_0_7_1_V(wire_ph_hit_o[0][7][1]),
.ph_hit_o_0_7_2_V(wire_ph_hit_o[0][7][2]),
.ph_hit_o_0_7_3_V(wire_ph_hit_o[0][7][3]),
.ph_hit_o_0_7_4_V(wire_ph_hit_o[0][7][4]),
.ph_hit_o_0_7_5_V(wire_ph_hit_o[0][7][5]),
.ph_hit_o_0_7_6_V(wire_ph_hit_o[0][7][6]),
.ph_hit_o_0_7_7_V(wire_ph_hit_o[0][7][7]),
.ph_hit_o_0_7_8_V(wire_ph_hit_o[0][7][8]),
.ph_hit_o_0_8_0_V(wire_ph_hit_o[0][8][0]),
.ph_hit_o_0_8_1_V(wire_ph_hit_o[0][8][1]),
.ph_hit_o_0_8_2_V(wire_ph_hit_o[0][8][2]),
.ph_hit_o_0_8_3_V(wire_ph_hit_o[0][8][3]),
.ph_hit_o_0_8_4_V(wire_ph_hit_o[0][8][4]),
.ph_hit_o_0_8_5_V(wire_ph_hit_o[0][8][5]),
.ph_hit_o_0_8_6_V(wire_ph_hit_o[0][8][6]),
.ph_hit_o_0_8_7_V(wire_ph_hit_o[0][8][7]),
.ph_hit_o_0_8_8_V(wire_ph_hit_o[0][8][8]),
.ph_hit_o_0_9_0_V(wire_ph_hit_o[0][9][0]),
.ph_hit_o_0_9_1_V(wire_ph_hit_o[0][9][1]),
.ph_hit_o_0_9_2_V(wire_ph_hit_o[0][9][2]),
.ph_hit_o_0_9_3_V(wire_ph_hit_o[0][9][3]),
.ph_hit_o_0_9_4_V(wire_ph_hit_o[0][9][4]),
.ph_hit_o_0_9_5_V(wire_ph_hit_o[0][9][5]),
.ph_hit_o_0_9_6_V(wire_ph_hit_o[0][9][6]),
.ph_hit_o_0_9_7_V(wire_ph_hit_o[0][9][7]),
.ph_hit_o_0_9_8_V(wire_ph_hit_o[0][9][8]),
.ph_hit_o_0_10_0_V(wire_ph_hit_o[0][10][0]),
.ph_hit_o_0_10_1_V(wire_ph_hit_o[0][10][1]),
.ph_hit_o_0_10_2_V(wire_ph_hit_o[0][10][2]),
.ph_hit_o_0_10_3_V(wire_ph_hit_o[0][10][3]),
.ph_hit_o_0_10_4_V(wire_ph_hit_o[0][10][4]),
.ph_hit_o_0_10_5_V(wire_ph_hit_o[0][10][5]),
.ph_hit_o_0_10_6_V(wire_ph_hit_o[0][10][6]),
.ph_hit_o_0_10_7_V(wire_ph_hit_o[0][10][7]),
.ph_hit_o_0_10_8_V(wire_ph_hit_o[0][10][8]),
.ph_hit_o_0_11_0_V(wire_ph_hit_o[0][11][0]),
.ph_hit_o_0_11_1_V(wire_ph_hit_o[0][11][1]),
.ph_hit_o_0_11_2_V(wire_ph_hit_o[0][11][2]),
.ph_hit_o_0_11_3_V(wire_ph_hit_o[0][11][3]),
.ph_hit_o_0_11_4_V(wire_ph_hit_o[0][11][4]),
.ph_hit_o_0_11_5_V(wire_ph_hit_o[0][11][5]),
.ph_hit_o_0_11_6_V(wire_ph_hit_o[0][11][6]),
.ph_hit_o_0_11_7_V(wire_ph_hit_o[0][11][7]),
.ph_hit_o_0_11_8_V(wire_ph_hit_o[0][11][8]),
.ph_hit_o_0_12_0_V(wire_ph_hit_o[0][12][0]),
.ph_hit_o_0_12_1_V(wire_ph_hit_o[0][12][1]),
.ph_hit_o_0_12_2_V(wire_ph_hit_o[0][12][2]),
.ph_hit_o_0_12_3_V(wire_ph_hit_o[0][12][3]),
.ph_hit_o_0_12_4_V(wire_ph_hit_o[0][12][4]),
.ph_hit_o_0_12_5_V(wire_ph_hit_o[0][12][5]),
.ph_hit_o_0_12_6_V(wire_ph_hit_o[0][12][6]),
.ph_hit_o_0_12_7_V(wire_ph_hit_o[0][12][7]),
.ph_hit_o_0_12_8_V(wire_ph_hit_o[0][12][8]),
.time_o_0_0_0_0_V_ap_vld(),
.time_o_0_0_0_1_V_ap_vld(),
.time_o_0_0_1_0_V_ap_vld(),
.time_o_0_0_1_1_V_ap_vld(),
.time_o_0_0_2_0_V_ap_vld(),
.time_o_0_0_2_1_V_ap_vld(),
.time_o_0_0_3_0_V_ap_vld(),
.time_o_0_0_3_1_V_ap_vld(),
.time_o_0_0_4_0_V_ap_vld(),
.time_o_0_0_4_1_V_ap_vld(),
.time_o_0_0_5_0_V_ap_vld(),
.time_o_0_0_5_1_V_ap_vld(),
.time_o_0_0_6_0_V_ap_vld(),
.time_o_0_0_6_1_V_ap_vld(),
.time_o_0_0_7_0_V_ap_vld(),
.time_o_0_0_7_1_V_ap_vld(),
.time_o_0_0_8_0_V_ap_vld(),
.time_o_0_0_8_1_V_ap_vld(),
.time_o_0_1_0_0_V_ap_vld(),
.time_o_0_1_0_1_V_ap_vld(),
.time_o_0_1_1_0_V_ap_vld(),
.time_o_0_1_1_1_V_ap_vld(),
.time_o_0_1_2_0_V_ap_vld(),
.time_o_0_1_2_1_V_ap_vld(),
.time_o_0_1_3_0_V_ap_vld(),
.time_o_0_1_3_1_V_ap_vld(),
.time_o_0_1_4_0_V_ap_vld(),
.time_o_0_1_4_1_V_ap_vld(),
.time_o_0_1_5_0_V_ap_vld(),
.time_o_0_1_5_1_V_ap_vld(),
.time_o_0_1_6_0_V_ap_vld(),
.time_o_0_1_6_1_V_ap_vld(),
.time_o_0_1_7_0_V_ap_vld(),
.time_o_0_1_7_1_V_ap_vld(),
.time_o_0_1_8_0_V_ap_vld(),
.time_o_0_1_8_1_V_ap_vld(),
.time_o_0_2_0_0_V_ap_vld(),
.time_o_0_2_0_1_V_ap_vld(),
.time_o_0_2_1_0_V_ap_vld(),
.time_o_0_2_1_1_V_ap_vld(),
.time_o_0_2_2_0_V_ap_vld(),
.time_o_0_2_2_1_V_ap_vld(),
.time_o_0_2_3_0_V_ap_vld(),
.time_o_0_2_3_1_V_ap_vld(),
.time_o_0_2_4_0_V_ap_vld(),
.time_o_0_2_4_1_V_ap_vld(),
.time_o_0_2_5_0_V_ap_vld(),
.time_o_0_2_5_1_V_ap_vld(),
.time_o_0_2_6_0_V_ap_vld(),
.time_o_0_2_6_1_V_ap_vld(),
.time_o_0_2_7_0_V_ap_vld(),
.time_o_0_2_7_1_V_ap_vld(),
.time_o_0_2_8_0_V_ap_vld(),
.time_o_0_2_8_1_V_ap_vld(),
.time_o_0_3_0_0_V_ap_vld(),
.time_o_0_3_0_1_V_ap_vld(),
.time_o_0_3_1_0_V_ap_vld(),
.time_o_0_3_1_1_V_ap_vld(),
.time_o_0_3_2_0_V_ap_vld(),
.time_o_0_3_2_1_V_ap_vld(),
.time_o_0_3_3_0_V_ap_vld(),
.time_o_0_3_3_1_V_ap_vld(),
.time_o_0_3_4_0_V_ap_vld(),
.time_o_0_3_4_1_V_ap_vld(),
.time_o_0_3_5_0_V_ap_vld(),
.time_o_0_3_5_1_V_ap_vld(),
.time_o_0_3_6_0_V_ap_vld(),
.time_o_0_3_6_1_V_ap_vld(),
.time_o_0_3_7_0_V_ap_vld(),
.time_o_0_3_7_1_V_ap_vld(),
.time_o_0_3_8_0_V_ap_vld(),
.time_o_0_3_8_1_V_ap_vld(),
.time_o_0_4_0_0_V_ap_vld(),
.time_o_0_4_0_1_V_ap_vld(),
.time_o_0_4_1_0_V_ap_vld(),
.time_o_0_4_1_1_V_ap_vld(),
.time_o_0_4_2_0_V_ap_vld(),
.time_o_0_4_2_1_V_ap_vld(),
.time_o_0_4_3_0_V_ap_vld(),
.time_o_0_4_3_1_V_ap_vld(),
.time_o_0_4_4_0_V_ap_vld(),
.time_o_0_4_4_1_V_ap_vld(),
.time_o_0_4_5_0_V_ap_vld(),
.time_o_0_4_5_1_V_ap_vld(),
.time_o_0_4_6_0_V_ap_vld(),
.time_o_0_4_6_1_V_ap_vld(),
.time_o_0_4_7_0_V_ap_vld(),
.time_o_0_4_7_1_V_ap_vld(),
.time_o_0_4_8_0_V_ap_vld(),
.time_o_0_4_8_1_V_ap_vld(),
.time_o_0_5_0_0_V_ap_vld(),
.time_o_0_5_0_1_V_ap_vld(),
.time_o_0_5_1_0_V_ap_vld(),
.time_o_0_5_1_1_V_ap_vld(),
.time_o_0_5_2_0_V_ap_vld(),
.time_o_0_5_2_1_V_ap_vld(),
.time_o_0_5_3_0_V_ap_vld(),
.time_o_0_5_3_1_V_ap_vld(),
.time_o_0_5_4_0_V_ap_vld(),
.time_o_0_5_4_1_V_ap_vld(),
.time_o_0_5_5_0_V_ap_vld(),
.time_o_0_5_5_1_V_ap_vld(),
.time_o_0_5_6_0_V_ap_vld(),
.time_o_0_5_6_1_V_ap_vld(),
.time_o_0_5_7_0_V_ap_vld(),
.time_o_0_5_7_1_V_ap_vld(),
.time_o_0_5_8_0_V_ap_vld(),
.time_o_0_5_8_1_V_ap_vld(),
.time_o_0_6_0_0_V_ap_vld(),
.time_o_0_6_0_1_V_ap_vld(),
.time_o_0_6_1_0_V_ap_vld(),
.time_o_0_6_1_1_V_ap_vld(),
.time_o_0_6_2_0_V_ap_vld(),
.time_o_0_6_2_1_V_ap_vld(),
.time_o_0_6_3_0_V_ap_vld(),
.time_o_0_6_3_1_V_ap_vld(),
.time_o_0_6_4_0_V_ap_vld(),
.time_o_0_6_4_1_V_ap_vld(),
.time_o_0_6_5_0_V_ap_vld(),
.time_o_0_6_5_1_V_ap_vld(),
.time_o_0_6_6_0_V_ap_vld(),
.time_o_0_6_6_1_V_ap_vld(),
.time_o_0_6_7_0_V_ap_vld(),
.time_o_0_6_7_1_V_ap_vld(),
.time_o_0_6_8_0_V_ap_vld(),
.time_o_0_6_8_1_V_ap_vld(),
.vl_o_0_0_0_V_ap_vld(),
.vl_o_0_0_1_V_ap_vld(),
.vl_o_0_0_2_V_ap_vld(),
.vl_o_0_0_3_V_ap_vld(),
.vl_o_0_0_4_V_ap_vld(),
.vl_o_0_0_5_V_ap_vld(),
.vl_o_0_0_6_V_ap_vld(),
.vl_o_0_0_7_V_ap_vld(),
.vl_o_0_0_8_V_ap_vld(),
.vl_o_0_1_0_V_ap_vld(),
.vl_o_0_1_1_V_ap_vld(),
.vl_o_0_1_2_V_ap_vld(),
.vl_o_0_1_3_V_ap_vld(),
.vl_o_0_1_4_V_ap_vld(),
.vl_o_0_1_5_V_ap_vld(),
.vl_o_0_1_6_V_ap_vld(),
.vl_o_0_1_7_V_ap_vld(),
.vl_o_0_1_8_V_ap_vld(),
.vl_o_0_2_0_V_ap_vld(),
.vl_o_0_2_1_V_ap_vld(),
.vl_o_0_2_2_V_ap_vld(),
.vl_o_0_2_3_V_ap_vld(),
.vl_o_0_2_4_V_ap_vld(),
.vl_o_0_2_5_V_ap_vld(),
.vl_o_0_2_6_V_ap_vld(),
.vl_o_0_2_7_V_ap_vld(),
.vl_o_0_2_8_V_ap_vld(),
.vl_o_0_3_0_V_ap_vld(),
.vl_o_0_3_1_V_ap_vld(),
.vl_o_0_3_2_V_ap_vld(),
.vl_o_0_3_3_V_ap_vld(),
.vl_o_0_3_4_V_ap_vld(),
.vl_o_0_3_5_V_ap_vld(),
.vl_o_0_3_6_V_ap_vld(),
.vl_o_0_3_7_V_ap_vld(),
.vl_o_0_3_8_V_ap_vld(),
.vl_o_0_4_0_V_ap_vld(),
.vl_o_0_4_1_V_ap_vld(),
.vl_o_0_4_2_V_ap_vld(),
.vl_o_0_4_3_V_ap_vld(),
.vl_o_0_4_4_V_ap_vld(),
.vl_o_0_4_5_V_ap_vld(),
.vl_o_0_4_6_V_ap_vld(),
.vl_o_0_4_7_V_ap_vld(),
.vl_o_0_4_8_V_ap_vld(),
.vl_o_0_5_0_V_ap_vld(),
.vl_o_0_5_1_V_ap_vld(),
.vl_o_0_5_2_V_ap_vld(),
.vl_o_0_5_3_V_ap_vld(),
.vl_o_0_5_4_V_ap_vld(),
.vl_o_0_5_5_V_ap_vld(),
.vl_o_0_5_6_V_ap_vld(),
.vl_o_0_5_7_V_ap_vld(),
.vl_o_0_5_8_V_ap_vld(),
.vl_o_0_6_0_V_ap_vld(),
.vl_o_0_6_1_V_ap_vld(),
.vl_o_0_6_2_V_ap_vld(),
.vl_o_0_6_3_V_ap_vld(),
.vl_o_0_6_4_V_ap_vld(),
.vl_o_0_6_5_V_ap_vld(),
.vl_o_0_6_6_V_ap_vld(),
.vl_o_0_6_7_V_ap_vld(),
.vl_o_0_6_8_V_ap_vld(),
.vl_o_0_7_0_V_ap_vld(),
.vl_o_0_7_1_V_ap_vld(),
.vl_o_0_7_2_V_ap_vld(),
.vl_o_0_7_3_V_ap_vld(),
.vl_o_0_7_4_V_ap_vld(),
.vl_o_0_7_5_V_ap_vld(),
.vl_o_0_7_6_V_ap_vld(),
.vl_o_0_7_7_V_ap_vld(),
.vl_o_0_7_8_V_ap_vld(),
.vl_o_0_8_0_V_ap_vld(),
.vl_o_0_8_1_V_ap_vld(),
.vl_o_0_8_2_V_ap_vld(),
.vl_o_0_8_3_V_ap_vld(),
.vl_o_0_8_4_V_ap_vld(),
.vl_o_0_8_5_V_ap_vld(),
.vl_o_0_8_6_V_ap_vld(),
.vl_o_0_8_7_V_ap_vld(),
.vl_o_0_8_8_V_ap_vld(),
.vl_o_0_9_0_V_ap_vld(),
.vl_o_0_9_1_V_ap_vld(),
.vl_o_0_9_2_V_ap_vld(),
.vl_o_0_9_3_V_ap_vld(),
.vl_o_0_9_4_V_ap_vld(),
.vl_o_0_9_5_V_ap_vld(),
.vl_o_0_9_6_V_ap_vld(),
.vl_o_0_9_7_V_ap_vld(),
.vl_o_0_9_8_V_ap_vld(),
.vl_o_0_10_0_V_ap_vld(),
.vl_o_0_10_1_V_ap_vld(),
.vl_o_0_10_2_V_ap_vld(),
.vl_o_0_10_3_V_ap_vld(),
.vl_o_0_10_4_V_ap_vld(),
.vl_o_0_10_5_V_ap_vld(),
.vl_o_0_10_6_V_ap_vld(),
.vl_o_0_10_7_V_ap_vld(),
.vl_o_0_10_8_V_ap_vld(),
.vl_o_0_11_0_V_ap_vld(),
.vl_o_0_11_1_V_ap_vld(),
.vl_o_0_11_2_V_ap_vld(),
.vl_o_0_11_3_V_ap_vld(),
.vl_o_0_11_4_V_ap_vld(),
.vl_o_0_11_5_V_ap_vld(),
.vl_o_0_11_6_V_ap_vld(),
.vl_o_0_11_7_V_ap_vld(),
.vl_o_0_11_8_V_ap_vld(),
.vl_o_0_12_0_V_ap_vld(),
.vl_o_0_12_1_V_ap_vld(),
.vl_o_0_12_2_V_ap_vld(),
.vl_o_0_12_3_V_ap_vld(),
.vl_o_0_12_4_V_ap_vld(),
.vl_o_0_12_5_V_ap_vld(),
.vl_o_0_12_6_V_ap_vld(),
.vl_o_0_12_7_V_ap_vld(),
.vl_o_0_12_8_V_ap_vld(),
.q_o_0_0_0_0_V_ap_vld(),
.q_o_0_0_0_1_V_ap_vld(),
.q_o_0_0_0_2_V_ap_vld(),
.q_o_0_0_1_0_V_ap_vld(),
.q_o_0_0_1_1_V_ap_vld(),
.q_o_0_0_1_2_V_ap_vld(),
.q_o_0_0_2_0_V_ap_vld(),
.q_o_0_0_2_1_V_ap_vld(),
.q_o_0_0_2_2_V_ap_vld(),
.q_o_0_0_3_0_V_ap_vld(),
.q_o_0_0_3_1_V_ap_vld(),
.q_o_0_0_3_2_V_ap_vld(),
.q_o_0_0_4_0_V_ap_vld(),
.q_o_0_0_4_1_V_ap_vld(),
.q_o_0_0_4_2_V_ap_vld(),
.q_o_0_0_5_0_V_ap_vld(),
.q_o_0_0_5_1_V_ap_vld(),
.q_o_0_0_5_2_V_ap_vld(),
.q_o_0_0_6_0_V_ap_vld(),
.q_o_0_0_6_1_V_ap_vld(),
.q_o_0_0_6_2_V_ap_vld(),
.q_o_0_0_7_0_V_ap_vld(),
.q_o_0_0_7_1_V_ap_vld(),
.q_o_0_0_7_2_V_ap_vld(),
.q_o_0_0_8_0_V_ap_vld(),
.q_o_0_0_8_1_V_ap_vld(),
.q_o_0_0_8_2_V_ap_vld(),
.q_o_0_1_0_0_V_ap_vld(),
.q_o_0_1_0_1_V_ap_vld(),
.q_o_0_1_0_2_V_ap_vld(),
.q_o_0_1_1_0_V_ap_vld(),
.q_o_0_1_1_1_V_ap_vld(),
.q_o_0_1_1_2_V_ap_vld(),
.q_o_0_1_2_0_V_ap_vld(),
.q_o_0_1_2_1_V_ap_vld(),
.q_o_0_1_2_2_V_ap_vld(),
.q_o_0_1_3_0_V_ap_vld(),
.q_o_0_1_3_1_V_ap_vld(),
.q_o_0_1_3_2_V_ap_vld(),
.q_o_0_1_4_0_V_ap_vld(),
.q_o_0_1_4_1_V_ap_vld(),
.q_o_0_1_4_2_V_ap_vld(),
.q_o_0_1_5_0_V_ap_vld(),
.q_o_0_1_5_1_V_ap_vld(),
.q_o_0_1_5_2_V_ap_vld(),
.q_o_0_1_6_0_V_ap_vld(),
.q_o_0_1_6_1_V_ap_vld(),
.q_o_0_1_6_2_V_ap_vld(),
.q_o_0_1_7_0_V_ap_vld(),
.q_o_0_1_7_1_V_ap_vld(),
.q_o_0_1_7_2_V_ap_vld(),
.q_o_0_1_8_0_V_ap_vld(),
.q_o_0_1_8_1_V_ap_vld(),
.q_o_0_1_8_2_V_ap_vld(),
.q_o_0_2_0_0_V_ap_vld(),
.q_o_0_2_0_1_V_ap_vld(),
.q_o_0_2_0_2_V_ap_vld(),
.q_o_0_2_1_0_V_ap_vld(),
.q_o_0_2_1_1_V_ap_vld(),
.q_o_0_2_1_2_V_ap_vld(),
.q_o_0_2_2_0_V_ap_vld(),
.q_o_0_2_2_1_V_ap_vld(),
.q_o_0_2_2_2_V_ap_vld(),
.q_o_0_2_3_0_V_ap_vld(),
.q_o_0_2_3_1_V_ap_vld(),
.q_o_0_2_3_2_V_ap_vld(),
.q_o_0_2_4_0_V_ap_vld(),
.q_o_0_2_4_1_V_ap_vld(),
.q_o_0_2_4_2_V_ap_vld(),
.q_o_0_2_5_0_V_ap_vld(),
.q_o_0_2_5_1_V_ap_vld(),
.q_o_0_2_5_2_V_ap_vld(),
.q_o_0_2_6_0_V_ap_vld(),
.q_o_0_2_6_1_V_ap_vld(),
.q_o_0_2_6_2_V_ap_vld(),
.q_o_0_2_7_0_V_ap_vld(),
.q_o_0_2_7_1_V_ap_vld(),
.q_o_0_2_7_2_V_ap_vld(),
.q_o_0_2_8_0_V_ap_vld(),
.q_o_0_2_8_1_V_ap_vld(),
.q_o_0_2_8_2_V_ap_vld(),
.q_o_0_3_0_0_V_ap_vld(),
.q_o_0_3_0_1_V_ap_vld(),
.q_o_0_3_0_2_V_ap_vld(),
.q_o_0_3_1_0_V_ap_vld(),
.q_o_0_3_1_1_V_ap_vld(),
.q_o_0_3_1_2_V_ap_vld(),
.q_o_0_3_2_0_V_ap_vld(),
.q_o_0_3_2_1_V_ap_vld(),
.q_o_0_3_2_2_V_ap_vld(),
.q_o_0_3_3_0_V_ap_vld(),
.q_o_0_3_3_1_V_ap_vld(),
.q_o_0_3_3_2_V_ap_vld(),
.q_o_0_3_4_0_V_ap_vld(),
.q_o_0_3_4_1_V_ap_vld(),
.q_o_0_3_4_2_V_ap_vld(),
.q_o_0_3_5_0_V_ap_vld(),
.q_o_0_3_5_1_V_ap_vld(),
.q_o_0_3_5_2_V_ap_vld(),
.q_o_0_3_6_0_V_ap_vld(),
.q_o_0_3_6_1_V_ap_vld(),
.q_o_0_3_6_2_V_ap_vld(),
.q_o_0_3_7_0_V_ap_vld(),
.q_o_0_3_7_1_V_ap_vld(),
.q_o_0_3_7_2_V_ap_vld(),
.q_o_0_3_8_0_V_ap_vld(),
.q_o_0_3_8_1_V_ap_vld(),
.q_o_0_3_8_2_V_ap_vld(),
.q_o_0_4_0_0_V_ap_vld(),
.q_o_0_4_0_1_V_ap_vld(),
.q_o_0_4_0_2_V_ap_vld(),
.q_o_0_4_1_0_V_ap_vld(),
.q_o_0_4_1_1_V_ap_vld(),
.q_o_0_4_1_2_V_ap_vld(),
.q_o_0_4_2_0_V_ap_vld(),
.q_o_0_4_2_1_V_ap_vld(),
.q_o_0_4_2_2_V_ap_vld(),
.q_o_0_4_3_0_V_ap_vld(),
.q_o_0_4_3_1_V_ap_vld(),
.q_o_0_4_3_2_V_ap_vld(),
.q_o_0_4_4_0_V_ap_vld(),
.q_o_0_4_4_1_V_ap_vld(),
.q_o_0_4_4_2_V_ap_vld(),
.q_o_0_4_5_0_V_ap_vld(),
.q_o_0_4_5_1_V_ap_vld(),
.q_o_0_4_5_2_V_ap_vld(),
.q_o_0_4_6_0_V_ap_vld(),
.q_o_0_4_6_1_V_ap_vld(),
.q_o_0_4_6_2_V_ap_vld(),
.q_o_0_4_7_0_V_ap_vld(),
.q_o_0_4_7_1_V_ap_vld(),
.q_o_0_4_7_2_V_ap_vld(),
.q_o_0_4_8_0_V_ap_vld(),
.q_o_0_4_8_1_V_ap_vld(),
.q_o_0_4_8_2_V_ap_vld(),
.q_o_0_5_0_0_V_ap_vld(),
.q_o_0_5_0_1_V_ap_vld(),
.q_o_0_5_0_2_V_ap_vld(),
.q_o_0_5_1_0_V_ap_vld(),
.q_o_0_5_1_1_V_ap_vld(),
.q_o_0_5_1_2_V_ap_vld(),
.q_o_0_5_2_0_V_ap_vld(),
.q_o_0_5_2_1_V_ap_vld(),
.q_o_0_5_2_2_V_ap_vld(),
.q_o_0_5_3_0_V_ap_vld(),
.q_o_0_5_3_1_V_ap_vld(),
.q_o_0_5_3_2_V_ap_vld(),
.q_o_0_5_4_0_V_ap_vld(),
.q_o_0_5_4_1_V_ap_vld(),
.q_o_0_5_4_2_V_ap_vld(),
.q_o_0_5_5_0_V_ap_vld(),
.q_o_0_5_5_1_V_ap_vld(),
.q_o_0_5_5_2_V_ap_vld(),
.q_o_0_5_6_0_V_ap_vld(),
.q_o_0_5_6_1_V_ap_vld(),
.q_o_0_5_6_2_V_ap_vld(),
.q_o_0_5_7_0_V_ap_vld(),
.q_o_0_5_7_1_V_ap_vld(),
.q_o_0_5_7_2_V_ap_vld(),
.q_o_0_5_8_0_V_ap_vld(),
.q_o_0_5_8_1_V_ap_vld(),
.q_o_0_5_8_2_V_ap_vld(),
.q_o_0_6_0_0_V_ap_vld(),
.q_o_0_6_0_1_V_ap_vld(),
.q_o_0_6_0_2_V_ap_vld(),
.q_o_0_6_1_0_V_ap_vld(),
.q_o_0_6_1_1_V_ap_vld(),
.q_o_0_6_1_2_V_ap_vld(),
.q_o_0_6_2_0_V_ap_vld(),
.q_o_0_6_2_1_V_ap_vld(),
.q_o_0_6_2_2_V_ap_vld(),
.q_o_0_6_3_0_V_ap_vld(),
.q_o_0_6_3_1_V_ap_vld(),
.q_o_0_6_3_2_V_ap_vld(),
.q_o_0_6_4_0_V_ap_vld(),
.q_o_0_6_4_1_V_ap_vld(),
.q_o_0_6_4_2_V_ap_vld(),
.q_o_0_6_5_0_V_ap_vld(),
.q_o_0_6_5_1_V_ap_vld(),
.q_o_0_6_5_2_V_ap_vld(),
.q_o_0_6_6_0_V_ap_vld(),
.q_o_0_6_6_1_V_ap_vld(),
.q_o_0_6_6_2_V_ap_vld(),
.q_o_0_6_7_0_V_ap_vld(),
.q_o_0_6_7_1_V_ap_vld(),
.q_o_0_6_7_2_V_ap_vld(),
.q_o_0_6_8_0_V_ap_vld(),
.q_o_0_6_8_1_V_ap_vld(),
.q_o_0_6_8_2_V_ap_vld(),
.q_o_0_7_0_0_V_ap_vld(),
.q_o_0_7_0_1_V_ap_vld(),
.q_o_0_7_0_2_V_ap_vld(),
.q_o_0_7_1_0_V_ap_vld(),
.q_o_0_7_1_1_V_ap_vld(),
.q_o_0_7_1_2_V_ap_vld(),
.q_o_0_7_2_0_V_ap_vld(),
.q_o_0_7_2_1_V_ap_vld(),
.q_o_0_7_2_2_V_ap_vld(),
.q_o_0_7_3_0_V_ap_vld(),
.q_o_0_7_3_1_V_ap_vld(),
.q_o_0_7_3_2_V_ap_vld(),
.q_o_0_7_4_0_V_ap_vld(),
.q_o_0_7_4_1_V_ap_vld(),
.q_o_0_7_4_2_V_ap_vld(),
.q_o_0_7_5_0_V_ap_vld(),
.q_o_0_7_5_1_V_ap_vld(),
.q_o_0_7_5_2_V_ap_vld(),
.q_o_0_7_6_0_V_ap_vld(),
.q_o_0_7_6_1_V_ap_vld(),
.q_o_0_7_6_2_V_ap_vld(),
.q_o_0_7_7_0_V_ap_vld(),
.q_o_0_7_7_1_V_ap_vld(),
.q_o_0_7_7_2_V_ap_vld(),
.q_o_0_7_8_0_V_ap_vld(),
.q_o_0_7_8_1_V_ap_vld(),
.q_o_0_7_8_2_V_ap_vld(),
.q_o_0_8_0_0_V_ap_vld(),
.q_o_0_8_0_1_V_ap_vld(),
.q_o_0_8_0_2_V_ap_vld(),
.q_o_0_8_1_0_V_ap_vld(),
.q_o_0_8_1_1_V_ap_vld(),
.q_o_0_8_1_2_V_ap_vld(),
.q_o_0_8_2_0_V_ap_vld(),
.q_o_0_8_2_1_V_ap_vld(),
.q_o_0_8_2_2_V_ap_vld(),
.q_o_0_8_3_0_V_ap_vld(),
.q_o_0_8_3_1_V_ap_vld(),
.q_o_0_8_3_2_V_ap_vld(),
.q_o_0_8_4_0_V_ap_vld(),
.q_o_0_8_4_1_V_ap_vld(),
.q_o_0_8_4_2_V_ap_vld(),
.q_o_0_8_5_0_V_ap_vld(),
.q_o_0_8_5_1_V_ap_vld(),
.q_o_0_8_5_2_V_ap_vld(),
.q_o_0_8_6_0_V_ap_vld(),
.q_o_0_8_6_1_V_ap_vld(),
.q_o_0_8_6_2_V_ap_vld(),
.q_o_0_8_7_0_V_ap_vld(),
.q_o_0_8_7_1_V_ap_vld(),
.q_o_0_8_7_2_V_ap_vld(),
.q_o_0_8_8_0_V_ap_vld(),
.q_o_0_8_8_1_V_ap_vld(),
.q_o_0_8_8_2_V_ap_vld(),
.q_o_0_9_0_0_V_ap_vld(),
.q_o_0_9_0_1_V_ap_vld(),
.q_o_0_9_0_2_V_ap_vld(),
.q_o_0_9_1_0_V_ap_vld(),
.q_o_0_9_1_1_V_ap_vld(),
.q_o_0_9_1_2_V_ap_vld(),
.q_o_0_9_2_0_V_ap_vld(),
.q_o_0_9_2_1_V_ap_vld(),
.q_o_0_9_2_2_V_ap_vld(),
.q_o_0_9_3_0_V_ap_vld(),
.q_o_0_9_3_1_V_ap_vld(),
.q_o_0_9_3_2_V_ap_vld(),
.q_o_0_9_4_0_V_ap_vld(),
.q_o_0_9_4_1_V_ap_vld(),
.q_o_0_9_4_2_V_ap_vld(),
.q_o_0_9_5_0_V_ap_vld(),
.q_o_0_9_5_1_V_ap_vld(),
.q_o_0_9_5_2_V_ap_vld(),
.q_o_0_9_6_0_V_ap_vld(),
.q_o_0_9_6_1_V_ap_vld(),
.q_o_0_9_6_2_V_ap_vld(),
.q_o_0_9_7_0_V_ap_vld(),
.q_o_0_9_7_1_V_ap_vld(),
.q_o_0_9_7_2_V_ap_vld(),
.q_o_0_9_8_0_V_ap_vld(),
.q_o_0_9_8_1_V_ap_vld(),
.q_o_0_9_8_2_V_ap_vld(),
.q_o_0_10_0_0_V_ap_vld(),
.q_o_0_10_0_1_V_ap_vld(),
.q_o_0_10_0_2_V_ap_vld(),
.q_o_0_10_1_0_V_ap_vld(),
.q_o_0_10_1_1_V_ap_vld(),
.q_o_0_10_1_2_V_ap_vld(),
.q_o_0_10_2_0_V_ap_vld(),
.q_o_0_10_2_1_V_ap_vld(),
.q_o_0_10_2_2_V_ap_vld(),
.q_o_0_10_3_0_V_ap_vld(),
.q_o_0_10_3_1_V_ap_vld(),
.q_o_0_10_3_2_V_ap_vld(),
.q_o_0_10_4_0_V_ap_vld(),
.q_o_0_10_4_1_V_ap_vld(),
.q_o_0_10_4_2_V_ap_vld(),
.q_o_0_10_5_0_V_ap_vld(),
.q_o_0_10_5_1_V_ap_vld(),
.q_o_0_10_5_2_V_ap_vld(),
.q_o_0_10_6_0_V_ap_vld(),
.q_o_0_10_6_1_V_ap_vld(),
.q_o_0_10_6_2_V_ap_vld(),
.q_o_0_10_7_0_V_ap_vld(),
.q_o_0_10_7_1_V_ap_vld(),
.q_o_0_10_7_2_V_ap_vld(),
.q_o_0_10_8_0_V_ap_vld(),
.q_o_0_10_8_1_V_ap_vld(),
.q_o_0_10_8_2_V_ap_vld(),
.q_o_0_11_0_0_V_ap_vld(),
.q_o_0_11_0_1_V_ap_vld(),
.q_o_0_11_0_2_V_ap_vld(),
.q_o_0_11_1_0_V_ap_vld(),
.q_o_0_11_1_1_V_ap_vld(),
.q_o_0_11_1_2_V_ap_vld(),
.q_o_0_11_2_0_V_ap_vld(),
.q_o_0_11_2_1_V_ap_vld(),
.q_o_0_11_2_2_V_ap_vld(),
.q_o_0_11_3_0_V_ap_vld(),
.q_o_0_11_3_1_V_ap_vld(),
.q_o_0_11_3_2_V_ap_vld(),
.q_o_0_11_4_0_V_ap_vld(),
.q_o_0_11_4_1_V_ap_vld(),
.q_o_0_11_4_2_V_ap_vld(),
.q_o_0_11_5_0_V_ap_vld(),
.q_o_0_11_5_1_V_ap_vld(),
.q_o_0_11_5_2_V_ap_vld(),
.q_o_0_11_6_0_V_ap_vld(),
.q_o_0_11_6_1_V_ap_vld(),
.q_o_0_11_6_2_V_ap_vld(),
.q_o_0_11_7_0_V_ap_vld(),
.q_o_0_11_7_1_V_ap_vld(),
.q_o_0_11_7_2_V_ap_vld(),
.q_o_0_11_8_0_V_ap_vld(),
.q_o_0_11_8_1_V_ap_vld(),
.q_o_0_11_8_2_V_ap_vld(),
.q_o_0_12_0_0_V_ap_vld(),
.q_o_0_12_0_1_V_ap_vld(),
.q_o_0_12_0_2_V_ap_vld(),
.q_o_0_12_1_0_V_ap_vld(),
.q_o_0_12_1_1_V_ap_vld(),
.q_o_0_12_1_2_V_ap_vld(),
.q_o_0_12_2_0_V_ap_vld(),
.q_o_0_12_2_1_V_ap_vld(),
.q_o_0_12_2_2_V_ap_vld(),
.q_o_0_12_3_0_V_ap_vld(),
.q_o_0_12_3_1_V_ap_vld(),
.q_o_0_12_3_2_V_ap_vld(),
.q_o_0_12_4_0_V_ap_vld(),
.q_o_0_12_4_1_V_ap_vld(),
.q_o_0_12_4_2_V_ap_vld(),
.q_o_0_12_5_0_V_ap_vld(),
.q_o_0_12_5_1_V_ap_vld(),
.q_o_0_12_5_2_V_ap_vld(),
.q_o_0_12_6_0_V_ap_vld(),
.q_o_0_12_6_1_V_ap_vld(),
.q_o_0_12_6_2_V_ap_vld(),
.q_o_0_12_7_0_V_ap_vld(),
.q_o_0_12_7_1_V_ap_vld(),
.q_o_0_12_7_2_V_ap_vld(),
.q_o_0_12_8_0_V_ap_vld(),
.q_o_0_12_8_1_V_ap_vld(),
.q_o_0_12_8_2_V_ap_vld(),
.cpatr_o_0_0_0_0_V_ap_vld(),
.cpatr_o_0_0_0_1_V_ap_vld(),
.cpatr_o_0_0_1_0_V_ap_vld(),
.cpatr_o_0_0_1_1_V_ap_vld(),
.cpatr_o_0_0_2_0_V_ap_vld(),
.cpatr_o_0_0_2_1_V_ap_vld(),
.cpatr_o_0_0_3_0_V_ap_vld(),
.cpatr_o_0_0_3_1_V_ap_vld(),
.cpatr_o_0_0_4_0_V_ap_vld(),
.cpatr_o_0_0_4_1_V_ap_vld(),
.cpatr_o_0_0_5_0_V_ap_vld(),
.cpatr_o_0_0_5_1_V_ap_vld(),
.cpatr_o_0_0_6_0_V_ap_vld(),
.cpatr_o_0_0_6_1_V_ap_vld(),
.cpatr_o_0_0_7_0_V_ap_vld(),
.cpatr_o_0_0_7_1_V_ap_vld(),
.cpatr_o_0_0_8_0_V_ap_vld(),
.cpatr_o_0_0_8_1_V_ap_vld(),
.cpatr_o_0_1_0_0_V_ap_vld(),
.cpatr_o_0_1_0_1_V_ap_vld(),
.cpatr_o_0_1_1_0_V_ap_vld(),
.cpatr_o_0_1_1_1_V_ap_vld(),
.cpatr_o_0_1_2_0_V_ap_vld(),
.cpatr_o_0_1_2_1_V_ap_vld(),
.cpatr_o_0_1_3_0_V_ap_vld(),
.cpatr_o_0_1_3_1_V_ap_vld(),
.cpatr_o_0_1_4_0_V_ap_vld(),
.cpatr_o_0_1_4_1_V_ap_vld(),
.cpatr_o_0_1_5_0_V_ap_vld(),
.cpatr_o_0_1_5_1_V_ap_vld(),
.cpatr_o_0_1_6_0_V_ap_vld(),
.cpatr_o_0_1_6_1_V_ap_vld(),
.cpatr_o_0_1_7_0_V_ap_vld(),
.cpatr_o_0_1_7_1_V_ap_vld(),
.cpatr_o_0_1_8_0_V_ap_vld(),
.cpatr_o_0_1_8_1_V_ap_vld(),
.cpatr_o_0_2_0_0_V_ap_vld(),
.cpatr_o_0_2_0_1_V_ap_vld(),
.cpatr_o_0_2_1_0_V_ap_vld(),
.cpatr_o_0_2_1_1_V_ap_vld(),
.cpatr_o_0_2_2_0_V_ap_vld(),
.cpatr_o_0_2_2_1_V_ap_vld(),
.cpatr_o_0_2_3_0_V_ap_vld(),
.cpatr_o_0_2_3_1_V_ap_vld(),
.cpatr_o_0_2_4_0_V_ap_vld(),
.cpatr_o_0_2_4_1_V_ap_vld(),
.cpatr_o_0_2_5_0_V_ap_vld(),
.cpatr_o_0_2_5_1_V_ap_vld(),
.cpatr_o_0_2_6_0_V_ap_vld(),
.cpatr_o_0_2_6_1_V_ap_vld(),
.cpatr_o_0_2_7_0_V_ap_vld(),
.cpatr_o_0_2_7_1_V_ap_vld(),
.cpatr_o_0_2_8_0_V_ap_vld(),
.cpatr_o_0_2_8_1_V_ap_vld(),
.cpatr_o_0_3_0_0_V_ap_vld(),
.cpatr_o_0_3_0_1_V_ap_vld(),
.cpatr_o_0_3_1_0_V_ap_vld(),
.cpatr_o_0_3_1_1_V_ap_vld(),
.cpatr_o_0_3_2_0_V_ap_vld(),
.cpatr_o_0_3_2_1_V_ap_vld(),
.cpatr_o_0_3_3_0_V_ap_vld(),
.cpatr_o_0_3_3_1_V_ap_vld(),
.cpatr_o_0_3_4_0_V_ap_vld(),
.cpatr_o_0_3_4_1_V_ap_vld(),
.cpatr_o_0_3_5_0_V_ap_vld(),
.cpatr_o_0_3_5_1_V_ap_vld(),
.cpatr_o_0_3_6_0_V_ap_vld(),
.cpatr_o_0_3_6_1_V_ap_vld(),
.cpatr_o_0_3_7_0_V_ap_vld(),
.cpatr_o_0_3_7_1_V_ap_vld(),
.cpatr_o_0_3_8_0_V_ap_vld(),
.cpatr_o_0_3_8_1_V_ap_vld(),
.cpatr_o_0_4_0_0_V_ap_vld(),
.cpatr_o_0_4_0_1_V_ap_vld(),
.cpatr_o_0_4_1_0_V_ap_vld(),
.cpatr_o_0_4_1_1_V_ap_vld(),
.cpatr_o_0_4_2_0_V_ap_vld(),
.cpatr_o_0_4_2_1_V_ap_vld(),
.cpatr_o_0_4_3_0_V_ap_vld(),
.cpatr_o_0_4_3_1_V_ap_vld(),
.cpatr_o_0_4_4_0_V_ap_vld(),
.cpatr_o_0_4_4_1_V_ap_vld(),
.cpatr_o_0_4_5_0_V_ap_vld(),
.cpatr_o_0_4_5_1_V_ap_vld(),
.cpatr_o_0_4_6_0_V_ap_vld(),
.cpatr_o_0_4_6_1_V_ap_vld(),
.cpatr_o_0_4_7_0_V_ap_vld(),
.cpatr_o_0_4_7_1_V_ap_vld(),
.cpatr_o_0_4_8_0_V_ap_vld(),
.cpatr_o_0_4_8_1_V_ap_vld(),
.cpatr_o_0_5_0_0_V_ap_vld(),
.cpatr_o_0_5_0_1_V_ap_vld(),
.cpatr_o_0_5_1_0_V_ap_vld(),
.cpatr_o_0_5_1_1_V_ap_vld(),
.cpatr_o_0_5_2_0_V_ap_vld(),
.cpatr_o_0_5_2_1_V_ap_vld(),
.cpatr_o_0_5_3_0_V_ap_vld(),
.cpatr_o_0_5_3_1_V_ap_vld(),
.cpatr_o_0_5_4_0_V_ap_vld(),
.cpatr_o_0_5_4_1_V_ap_vld(),
.cpatr_o_0_5_5_0_V_ap_vld(),
.cpatr_o_0_5_5_1_V_ap_vld(),
.cpatr_o_0_5_6_0_V_ap_vld(),
.cpatr_o_0_5_6_1_V_ap_vld(),
.cpatr_o_0_5_7_0_V_ap_vld(),
.cpatr_o_0_5_7_1_V_ap_vld(),
.cpatr_o_0_5_8_0_V_ap_vld(),
.cpatr_o_0_5_8_1_V_ap_vld(),
.ph_o_0_0_0_0_V_ap_vld(),
.ph_o_0_0_0_1_V_ap_vld(),
.ph_o_0_0_1_0_V_ap_vld(),
.ph_o_0_0_1_1_V_ap_vld(),
.ph_o_0_0_2_0_V_ap_vld(),
.ph_o_0_0_2_1_V_ap_vld(),
.ph_o_0_0_3_0_V_ap_vld(),
.ph_o_0_0_3_1_V_ap_vld(),
.ph_o_0_0_4_0_V_ap_vld(),
.ph_o_0_0_4_1_V_ap_vld(),
.ph_o_0_0_5_0_V_ap_vld(),
.ph_o_0_0_5_1_V_ap_vld(),
.ph_o_0_0_6_0_V_ap_vld(),
.ph_o_0_0_6_1_V_ap_vld(),
.ph_o_0_0_7_0_V_ap_vld(),
.ph_o_0_0_7_1_V_ap_vld(),
.ph_o_0_0_8_0_V_ap_vld(),
.ph_o_0_0_8_1_V_ap_vld(),
.ph_o_0_1_0_0_V_ap_vld(),
.ph_o_0_1_0_1_V_ap_vld(),
.ph_o_0_1_1_0_V_ap_vld(),
.ph_o_0_1_1_1_V_ap_vld(),
.ph_o_0_1_2_0_V_ap_vld(),
.ph_o_0_1_2_1_V_ap_vld(),
.ph_o_0_1_3_0_V_ap_vld(),
.ph_o_0_1_3_1_V_ap_vld(),
.ph_o_0_1_4_0_V_ap_vld(),
.ph_o_0_1_4_1_V_ap_vld(),
.ph_o_0_1_5_0_V_ap_vld(),
.ph_o_0_1_5_1_V_ap_vld(),
.ph_o_0_1_6_0_V_ap_vld(),
.ph_o_0_1_6_1_V_ap_vld(),
.ph_o_0_1_7_0_V_ap_vld(),
.ph_o_0_1_7_1_V_ap_vld(),
.ph_o_0_1_8_0_V_ap_vld(),
.ph_o_0_1_8_1_V_ap_vld(),
.ph_o_0_2_0_0_V_ap_vld(),
.ph_o_0_2_0_1_V_ap_vld(),
.ph_o_0_2_1_0_V_ap_vld(),
.ph_o_0_2_1_1_V_ap_vld(),
.ph_o_0_2_2_0_V_ap_vld(),
.ph_o_0_2_2_1_V_ap_vld(),
.ph_o_0_2_3_0_V_ap_vld(),
.ph_o_0_2_3_1_V_ap_vld(),
.ph_o_0_2_4_0_V_ap_vld(),
.ph_o_0_2_4_1_V_ap_vld(),
.ph_o_0_2_5_0_V_ap_vld(),
.ph_o_0_2_5_1_V_ap_vld(),
.ph_o_0_2_6_0_V_ap_vld(),
.ph_o_0_2_6_1_V_ap_vld(),
.ph_o_0_2_7_0_V_ap_vld(),
.ph_o_0_2_7_1_V_ap_vld(),
.ph_o_0_2_8_0_V_ap_vld(),
.ph_o_0_2_8_1_V_ap_vld(),
.ph_o_0_3_0_0_V_ap_vld(),
.ph_o_0_3_0_1_V_ap_vld(),
.ph_o_0_3_1_0_V_ap_vld(),
.ph_o_0_3_1_1_V_ap_vld(),
.ph_o_0_3_2_0_V_ap_vld(),
.ph_o_0_3_2_1_V_ap_vld(),
.ph_o_0_3_3_0_V_ap_vld(),
.ph_o_0_3_3_1_V_ap_vld(),
.ph_o_0_3_4_0_V_ap_vld(),
.ph_o_0_3_4_1_V_ap_vld(),
.ph_o_0_3_5_0_V_ap_vld(),
.ph_o_0_3_5_1_V_ap_vld(),
.ph_o_0_3_6_0_V_ap_vld(),
.ph_o_0_3_6_1_V_ap_vld(),
.ph_o_0_3_7_0_V_ap_vld(),
.ph_o_0_3_7_1_V_ap_vld(),
.ph_o_0_3_8_0_V_ap_vld(),
.ph_o_0_3_8_1_V_ap_vld(),
.ph_o_0_4_0_0_V_ap_vld(),
.ph_o_0_4_0_1_V_ap_vld(),
.ph_o_0_4_1_0_V_ap_vld(),
.ph_o_0_4_1_1_V_ap_vld(),
.ph_o_0_4_2_0_V_ap_vld(),
.ph_o_0_4_2_1_V_ap_vld(),
.ph_o_0_4_3_0_V_ap_vld(),
.ph_o_0_4_3_1_V_ap_vld(),
.ph_o_0_4_4_0_V_ap_vld(),
.ph_o_0_4_4_1_V_ap_vld(),
.ph_o_0_4_5_0_V_ap_vld(),
.ph_o_0_4_5_1_V_ap_vld(),
.ph_o_0_4_6_0_V_ap_vld(),
.ph_o_0_4_6_1_V_ap_vld(),
.ph_o_0_4_7_0_V_ap_vld(),
.ph_o_0_4_7_1_V_ap_vld(),
.ph_o_0_4_8_0_V_ap_vld(),
.ph_o_0_4_8_1_V_ap_vld(),
.ph_o_0_5_0_0_V_ap_vld(),
.ph_o_0_5_0_1_V_ap_vld(),
.ph_o_0_5_1_0_V_ap_vld(),
.ph_o_0_5_1_1_V_ap_vld(),
.ph_o_0_5_2_0_V_ap_vld(),
.ph_o_0_5_2_1_V_ap_vld(),
.ph_o_0_5_3_0_V_ap_vld(),
.ph_o_0_5_3_1_V_ap_vld(),
.ph_o_0_5_4_0_V_ap_vld(),
.ph_o_0_5_4_1_V_ap_vld(),
.ph_o_0_5_5_0_V_ap_vld(),
.ph_o_0_5_5_1_V_ap_vld(),
.ph_o_0_5_6_0_V_ap_vld(),
.ph_o_0_5_6_1_V_ap_vld(),
.ph_o_0_5_7_0_V_ap_vld(),
.ph_o_0_5_7_1_V_ap_vld(),
.ph_o_0_5_8_0_V_ap_vld(),
.ph_o_0_5_8_1_V_ap_vld(),
.th11_o_0_0_0_0_V_ap_vld(),
.th11_o_0_0_0_1_V_ap_vld(),
.th11_o_0_0_1_0_V_ap_vld(),
.th11_o_0_0_1_1_V_ap_vld(),
.th11_o_0_0_2_0_V_ap_vld(),
.th11_o_0_0_2_1_V_ap_vld(),
.th11_o_0_0_3_0_V_ap_vld(),
.th11_o_0_0_3_1_V_ap_vld(),
.th11_o_0_0_4_0_V_ap_vld(),
.th11_o_0_0_4_1_V_ap_vld(),
.th11_o_0_0_5_0_V_ap_vld(),
.th11_o_0_0_5_1_V_ap_vld(),
.th11_o_0_0_6_0_V_ap_vld(),
.th11_o_0_0_6_1_V_ap_vld(),
.th11_o_0_0_7_0_V_ap_vld(),
.th11_o_0_0_7_1_V_ap_vld(),
.th11_o_0_0_8_0_V_ap_vld(),
.th11_o_0_0_8_1_V_ap_vld(),
.th11_o_0_1_0_0_V_ap_vld(),
.th11_o_0_1_0_1_V_ap_vld(),
.th11_o_0_1_1_0_V_ap_vld(),
.th11_o_0_1_1_1_V_ap_vld(),
.th11_o_0_1_2_0_V_ap_vld(),
.th11_o_0_1_2_1_V_ap_vld(),
.th11_o_0_1_3_0_V_ap_vld(),
.th11_o_0_1_3_1_V_ap_vld(),
.th11_o_0_1_4_0_V_ap_vld(),
.th11_o_0_1_4_1_V_ap_vld(),
.th11_o_0_1_5_0_V_ap_vld(),
.th11_o_0_1_5_1_V_ap_vld(),
.th11_o_0_1_6_0_V_ap_vld(),
.th11_o_0_1_6_1_V_ap_vld(),
.th11_o_0_1_7_0_V_ap_vld(),
.th11_o_0_1_7_1_V_ap_vld(),
.th11_o_0_1_8_0_V_ap_vld(),
.th11_o_0_1_8_1_V_ap_vld(),
.th11_o_0_2_0_0_V_ap_vld(),
.th11_o_0_2_0_1_V_ap_vld(),
.th11_o_0_2_1_0_V_ap_vld(),
.th11_o_0_2_1_1_V_ap_vld(),
.th11_o_0_2_2_0_V_ap_vld(),
.th11_o_0_2_2_1_V_ap_vld(),
.th11_o_0_2_3_0_V_ap_vld(),
.th11_o_0_2_3_1_V_ap_vld(),
.th11_o_0_2_4_0_V_ap_vld(),
.th11_o_0_2_4_1_V_ap_vld(),
.th11_o_0_2_5_0_V_ap_vld(),
.th11_o_0_2_5_1_V_ap_vld(),
.th11_o_0_2_6_0_V_ap_vld(),
.th11_o_0_2_6_1_V_ap_vld(),
.th11_o_0_2_7_0_V_ap_vld(),
.th11_o_0_2_7_1_V_ap_vld(),
.th11_o_0_2_8_0_V_ap_vld(),
.th11_o_0_2_8_1_V_ap_vld(),
.th11_o_0_3_0_0_V_ap_vld(),
.th11_o_0_3_0_1_V_ap_vld(),
.th11_o_0_3_1_0_V_ap_vld(),
.th11_o_0_3_1_1_V_ap_vld(),
.th11_o_0_3_2_0_V_ap_vld(),
.th11_o_0_3_2_1_V_ap_vld(),
.th11_o_0_3_3_0_V_ap_vld(),
.th11_o_0_3_3_1_V_ap_vld(),
.th11_o_0_3_4_0_V_ap_vld(),
.th11_o_0_3_4_1_V_ap_vld(),
.th11_o_0_3_5_0_V_ap_vld(),
.th11_o_0_3_5_1_V_ap_vld(),
.th11_o_0_3_6_0_V_ap_vld(),
.th11_o_0_3_6_1_V_ap_vld(),
.th11_o_0_3_7_0_V_ap_vld(),
.th11_o_0_3_7_1_V_ap_vld(),
.th11_o_0_3_8_0_V_ap_vld(),
.th11_o_0_3_8_1_V_ap_vld(),
.th11_o_0_4_0_0_V_ap_vld(),
.th11_o_0_4_0_1_V_ap_vld(),
.th11_o_0_4_1_0_V_ap_vld(),
.th11_o_0_4_1_1_V_ap_vld(),
.th11_o_0_4_2_0_V_ap_vld(),
.th11_o_0_4_2_1_V_ap_vld(),
.th11_o_0_4_3_0_V_ap_vld(),
.th11_o_0_4_3_1_V_ap_vld(),
.th11_o_0_4_4_0_V_ap_vld(),
.th11_o_0_4_4_1_V_ap_vld(),
.th11_o_0_4_5_0_V_ap_vld(),
.th11_o_0_4_5_1_V_ap_vld(),
.th11_o_0_4_6_0_V_ap_vld(),
.th11_o_0_4_6_1_V_ap_vld(),
.th11_o_0_4_7_0_V_ap_vld(),
.th11_o_0_4_7_1_V_ap_vld(),
.th11_o_0_4_8_0_V_ap_vld(),
.th11_o_0_4_8_1_V_ap_vld(),
.th11_o_0_5_0_0_V_ap_vld(),
.th11_o_0_5_0_1_V_ap_vld(),
.th11_o_0_5_1_0_V_ap_vld(),
.th11_o_0_5_1_1_V_ap_vld(),
.th11_o_0_5_2_0_V_ap_vld(),
.th11_o_0_5_2_1_V_ap_vld(),
.th11_o_0_5_3_0_V_ap_vld(),
.th11_o_0_5_3_1_V_ap_vld(),
.th11_o_0_5_4_0_V_ap_vld(),
.th11_o_0_5_4_1_V_ap_vld(),
.th11_o_0_5_5_0_V_ap_vld(),
.th11_o_0_5_5_1_V_ap_vld(),
.th11_o_0_5_6_0_V_ap_vld(),
.th11_o_0_5_6_1_V_ap_vld(),
.th11_o_0_5_7_0_V_ap_vld(),
.th11_o_0_5_7_1_V_ap_vld(),
.th11_o_0_5_8_0_V_ap_vld(),
.th11_o_0_5_8_1_V_ap_vld(),
.th_o_0_0_0_0_V_ap_vld(),
.th_o_0_0_0_1_V_ap_vld(),
.th_o_0_0_0_2_V_ap_vld(),
.th_o_0_0_0_3_V_ap_vld(),
.th_o_0_0_1_0_V_ap_vld(),
.th_o_0_0_1_1_V_ap_vld(),
.th_o_0_0_1_2_V_ap_vld(),
.th_o_0_0_1_3_V_ap_vld(),
.th_o_0_0_2_0_V_ap_vld(),
.th_o_0_0_2_1_V_ap_vld(),
.th_o_0_0_2_2_V_ap_vld(),
.th_o_0_0_2_3_V_ap_vld(),
.th_o_0_1_0_0_V_ap_vld(),
.th_o_0_1_0_1_V_ap_vld(),
.th_o_0_1_0_2_V_ap_vld(),
.th_o_0_1_0_3_V_ap_vld(),
.th_o_0_1_1_0_V_ap_vld(),
.th_o_0_1_1_1_V_ap_vld(),
.th_o_0_1_1_2_V_ap_vld(),
.th_o_0_1_1_3_V_ap_vld(),
.th_o_0_1_2_0_V_ap_vld(),
.th_o_0_1_2_1_V_ap_vld(),
.th_o_0_1_2_2_V_ap_vld(),
.th_o_0_1_2_3_V_ap_vld(),
.th_o_0_2_0_0_V_ap_vld(),
.th_o_0_2_0_1_V_ap_vld(),
.th_o_0_2_0_2_V_ap_vld(),
.th_o_0_2_0_3_V_ap_vld(),
.th_o_0_2_1_0_V_ap_vld(),
.th_o_0_2_1_1_V_ap_vld(),
.th_o_0_2_1_2_V_ap_vld(),
.th_o_0_2_1_3_V_ap_vld(),
.th_o_0_2_2_0_V_ap_vld(),
.th_o_0_2_2_1_V_ap_vld(),
.th_o_0_2_2_2_V_ap_vld(),
.th_o_0_2_2_3_V_ap_vld(),
.phzvl_o_0_0_0_V_ap_vld(),
.phzvl_o_0_0_1_V_ap_vld(),
.phzvl_o_0_0_2_V_ap_vld(),
.phzvl_o_0_0_3_V_ap_vld(),
.phzvl_o_0_0_4_V_ap_vld(),
.phzvl_o_0_0_5_V_ap_vld(),
.phzvl_o_0_0_6_V_ap_vld(),
.phzvl_o_0_0_7_V_ap_vld(),
.phzvl_o_0_0_8_V_ap_vld(),
.phzvl_o_0_1_0_V_ap_vld(),
.phzvl_o_0_1_1_V_ap_vld(),
.phzvl_o_0_1_2_V_ap_vld(),
.phzvl_o_0_1_3_V_ap_vld(),
.phzvl_o_0_1_4_V_ap_vld(),
.phzvl_o_0_1_5_V_ap_vld(),
.phzvl_o_0_1_6_V_ap_vld(),
.phzvl_o_0_1_7_V_ap_vld(),
.phzvl_o_0_1_8_V_ap_vld(),
.phzvl_o_0_2_0_V_ap_vld(),
.phzvl_o_0_2_1_V_ap_vld(),
.phzvl_o_0_2_2_V_ap_vld(),
.phzvl_o_0_2_3_V_ap_vld(),
.phzvl_o_0_2_4_V_ap_vld(),
.phzvl_o_0_2_5_V_ap_vld(),
.phzvl_o_0_2_6_V_ap_vld(),
.phzvl_o_0_2_7_V_ap_vld(),
.phzvl_o_0_2_8_V_ap_vld(),
.phzvl_o_0_3_0_V_ap_vld(),
.phzvl_o_0_3_1_V_ap_vld(),
.phzvl_o_0_3_2_V_ap_vld(),
.phzvl_o_0_3_3_V_ap_vld(),
.phzvl_o_0_3_4_V_ap_vld(),
.phzvl_o_0_3_5_V_ap_vld(),
.phzvl_o_0_3_6_V_ap_vld(),
.phzvl_o_0_3_7_V_ap_vld(),
.phzvl_o_0_3_8_V_ap_vld(),
.phzvl_o_0_4_0_V_ap_vld(),
.phzvl_o_0_4_1_V_ap_vld(),
.phzvl_o_0_4_2_V_ap_vld(),
.phzvl_o_0_4_3_V_ap_vld(),
.phzvl_o_0_4_4_V_ap_vld(),
.phzvl_o_0_4_5_V_ap_vld(),
.phzvl_o_0_4_6_V_ap_vld(),
.phzvl_o_0_4_7_V_ap_vld(),
.phzvl_o_0_4_8_V_ap_vld(),
.phzvl_o_0_5_0_V_ap_vld(),
.phzvl_o_0_5_1_V_ap_vld(),
.phzvl_o_0_5_2_V_ap_vld(),
.phzvl_o_0_5_3_V_ap_vld(),
.phzvl_o_0_5_4_V_ap_vld(),
.phzvl_o_0_5_5_V_ap_vld(),
.phzvl_o_0_5_6_V_ap_vld(),
.phzvl_o_0_5_7_V_ap_vld(),
.phzvl_o_0_5_8_V_ap_vld(),
.phzvl_o_0_6_0_V_ap_vld(),
.phzvl_o_0_6_1_V_ap_vld(),
.phzvl_o_0_6_2_V_ap_vld(),
.phzvl_o_0_6_3_V_ap_vld(),
.phzvl_o_0_6_4_V_ap_vld(),
.phzvl_o_0_6_5_V_ap_vld(),
.phzvl_o_0_6_6_V_ap_vld(),
.phzvl_o_0_6_7_V_ap_vld(),
.phzvl_o_0_6_8_V_ap_vld(),
.phzvl_o_0_7_0_V_ap_vld(),
.phzvl_o_0_7_1_V_ap_vld(),
.phzvl_o_0_7_2_V_ap_vld(),
.phzvl_o_0_7_3_V_ap_vld(),
.phzvl_o_0_7_4_V_ap_vld(),
.phzvl_o_0_7_5_V_ap_vld(),
.phzvl_o_0_7_6_V_ap_vld(),
.phzvl_o_0_7_7_V_ap_vld(),
.phzvl_o_0_7_8_V_ap_vld(),
.phzvl_o_0_8_0_V_ap_vld(),
.phzvl_o_0_8_1_V_ap_vld(),
.phzvl_o_0_8_2_V_ap_vld(),
.phzvl_o_0_8_3_V_ap_vld(),
.phzvl_o_0_8_4_V_ap_vld(),
.phzvl_o_0_8_5_V_ap_vld(),
.phzvl_o_0_8_6_V_ap_vld(),
.phzvl_o_0_8_7_V_ap_vld(),
.phzvl_o_0_8_8_V_ap_vld(),
.phzvl_o_0_9_0_V_ap_vld(),
.phzvl_o_0_9_1_V_ap_vld(),
.phzvl_o_0_9_2_V_ap_vld(),
.phzvl_o_0_9_3_V_ap_vld(),
.phzvl_o_0_9_4_V_ap_vld(),
.phzvl_o_0_9_5_V_ap_vld(),
.phzvl_o_0_9_6_V_ap_vld(),
.phzvl_o_0_9_7_V_ap_vld(),
.phzvl_o_0_9_8_V_ap_vld(),
.phzvl_o_0_10_0_V_ap_vld(),
.phzvl_o_0_10_1_V_ap_vld(),
.phzvl_o_0_10_2_V_ap_vld(),
.phzvl_o_0_10_3_V_ap_vld(),
.phzvl_o_0_10_4_V_ap_vld(),
.phzvl_o_0_10_5_V_ap_vld(),
.phzvl_o_0_10_6_V_ap_vld(),
.phzvl_o_0_10_7_V_ap_vld(),
.phzvl_o_0_10_8_V_ap_vld(),
.phzvl_o_0_11_0_V_ap_vld(),
.phzvl_o_0_11_1_V_ap_vld(),
.phzvl_o_0_11_2_V_ap_vld(),
.phzvl_o_0_11_3_V_ap_vld(),
.phzvl_o_0_11_4_V_ap_vld(),
.phzvl_o_0_11_5_V_ap_vld(),
.phzvl_o_0_11_6_V_ap_vld(),
.phzvl_o_0_11_7_V_ap_vld(),
.phzvl_o_0_11_8_V_ap_vld(),
.phzvl_o_0_12_0_V_ap_vld(),
.phzvl_o_0_12_1_V_ap_vld(),
.phzvl_o_0_12_2_V_ap_vld(),
.phzvl_o_0_12_3_V_ap_vld(),
.phzvl_o_0_12_4_V_ap_vld(),
.phzvl_o_0_12_5_V_ap_vld(),
.phzvl_o_0_12_6_V_ap_vld(),
.phzvl_o_0_12_7_V_ap_vld(),
.phzvl_o_0_12_8_V_ap_vld(),
.ph_hit_o_0_0_0_V_ap_vld(),
.ph_hit_o_0_0_1_V_ap_vld(),
.ph_hit_o_0_0_2_V_ap_vld(),
.ph_hit_o_0_0_3_V_ap_vld(),
.ph_hit_o_0_0_4_V_ap_vld(),
.ph_hit_o_0_0_5_V_ap_vld(),
.ph_hit_o_0_0_6_V_ap_vld(),
.ph_hit_o_0_0_7_V_ap_vld(),
.ph_hit_o_0_0_8_V_ap_vld(),
.ph_hit_o_0_1_0_V_ap_vld(),
.ph_hit_o_0_1_1_V_ap_vld(),
.ph_hit_o_0_1_2_V_ap_vld(),
.ph_hit_o_0_1_3_V_ap_vld(),
.ph_hit_o_0_1_4_V_ap_vld(),
.ph_hit_o_0_1_5_V_ap_vld(),
.ph_hit_o_0_1_6_V_ap_vld(),
.ph_hit_o_0_1_7_V_ap_vld(),
.ph_hit_o_0_1_8_V_ap_vld(),
.ph_hit_o_0_2_0_V_ap_vld(),
.ph_hit_o_0_2_1_V_ap_vld(),
.ph_hit_o_0_2_2_V_ap_vld(),
.ph_hit_o_0_2_3_V_ap_vld(),
.ph_hit_o_0_2_4_V_ap_vld(),
.ph_hit_o_0_2_5_V_ap_vld(),
.ph_hit_o_0_2_6_V_ap_vld(),
.ph_hit_o_0_2_7_V_ap_vld(),
.ph_hit_o_0_2_8_V_ap_vld(),
.ph_hit_o_0_3_0_V_ap_vld(),
.ph_hit_o_0_3_1_V_ap_vld(),
.ph_hit_o_0_3_2_V_ap_vld(),
.ph_hit_o_0_3_3_V_ap_vld(),
.ph_hit_o_0_3_4_V_ap_vld(),
.ph_hit_o_0_3_5_V_ap_vld(),
.ph_hit_o_0_3_6_V_ap_vld(),
.ph_hit_o_0_3_7_V_ap_vld(),
.ph_hit_o_0_3_8_V_ap_vld(),
.ph_hit_o_0_4_0_V_ap_vld(),
.ph_hit_o_0_4_1_V_ap_vld(),
.ph_hit_o_0_4_2_V_ap_vld(),
.ph_hit_o_0_4_3_V_ap_vld(),
.ph_hit_o_0_4_4_V_ap_vld(),
.ph_hit_o_0_4_5_V_ap_vld(),
.ph_hit_o_0_4_6_V_ap_vld(),
.ph_hit_o_0_4_7_V_ap_vld(),
.ph_hit_o_0_4_8_V_ap_vld(),
.ph_hit_o_0_5_0_V_ap_vld(),
.ph_hit_o_0_5_1_V_ap_vld(),
.ph_hit_o_0_5_2_V_ap_vld(),
.ph_hit_o_0_5_3_V_ap_vld(),
.ph_hit_o_0_5_4_V_ap_vld(),
.ph_hit_o_0_5_5_V_ap_vld(),
.ph_hit_o_0_5_6_V_ap_vld(),
.ph_hit_o_0_5_7_V_ap_vld(),
.ph_hit_o_0_5_8_V_ap_vld(),
.ph_hit_o_0_6_0_V_ap_vld(),
.ph_hit_o_0_6_1_V_ap_vld(),
.ph_hit_o_0_6_2_V_ap_vld(),
.ph_hit_o_0_6_3_V_ap_vld(),
.ph_hit_o_0_6_4_V_ap_vld(),
.ph_hit_o_0_6_5_V_ap_vld(),
.ph_hit_o_0_6_6_V_ap_vld(),
.ph_hit_o_0_6_7_V_ap_vld(),
.ph_hit_o_0_6_8_V_ap_vld(),
.ph_hit_o_0_7_0_V_ap_vld(),
.ph_hit_o_0_7_1_V_ap_vld(),
.ph_hit_o_0_7_2_V_ap_vld(),
.ph_hit_o_0_7_3_V_ap_vld(),
.ph_hit_o_0_7_4_V_ap_vld(),
.ph_hit_o_0_7_5_V_ap_vld(),
.ph_hit_o_0_7_6_V_ap_vld(),
.ph_hit_o_0_7_7_V_ap_vld(),
.ph_hit_o_0_7_8_V_ap_vld(),
.ph_hit_o_0_8_0_V_ap_vld(),
.ph_hit_o_0_8_1_V_ap_vld(),
.ph_hit_o_0_8_2_V_ap_vld(),
.ph_hit_o_0_8_3_V_ap_vld(),
.ph_hit_o_0_8_4_V_ap_vld(),
.ph_hit_o_0_8_5_V_ap_vld(),
.ph_hit_o_0_8_6_V_ap_vld(),
.ph_hit_o_0_8_7_V_ap_vld(),
.ph_hit_o_0_8_8_V_ap_vld(),
.ph_hit_o_0_9_0_V_ap_vld(),
.ph_hit_o_0_9_1_V_ap_vld(),
.ph_hit_o_0_9_2_V_ap_vld(),
.ph_hit_o_0_9_3_V_ap_vld(),
.ph_hit_o_0_9_4_V_ap_vld(),
.ph_hit_o_0_9_5_V_ap_vld(),
.ph_hit_o_0_9_6_V_ap_vld(),
.ph_hit_o_0_9_7_V_ap_vld(),
.ph_hit_o_0_9_8_V_ap_vld(),
.ph_hit_o_0_10_0_V_ap_vld(),
.ph_hit_o_0_10_1_V_ap_vld(),
.ph_hit_o_0_10_2_V_ap_vld(),
.ph_hit_o_0_10_3_V_ap_vld(),
.ph_hit_o_0_10_4_V_ap_vld(),
.ph_hit_o_0_10_5_V_ap_vld(),
.ph_hit_o_0_10_6_V_ap_vld(),
.ph_hit_o_0_10_7_V_ap_vld(),
.ph_hit_o_0_10_8_V_ap_vld(),
.ph_hit_o_0_11_0_V_ap_vld(),
.ph_hit_o_0_11_1_V_ap_vld(),
.ph_hit_o_0_11_2_V_ap_vld(),
.ph_hit_o_0_11_3_V_ap_vld(),
.ph_hit_o_0_11_4_V_ap_vld(),
.ph_hit_o_0_11_5_V_ap_vld(),
.ph_hit_o_0_11_6_V_ap_vld(),
.ph_hit_o_0_11_7_V_ap_vld(),
.ph_hit_o_0_11_8_V_ap_vld(),
.ph_hit_o_0_12_0_V_ap_vld(),
.ph_hit_o_0_12_1_V_ap_vld(),
.ph_hit_o_0_12_2_V_ap_vld(),
.ph_hit_o_0_12_3_V_ap_vld(),
.ph_hit_o_0_12_4_V_ap_vld(),
.ph_hit_o_0_12_5_V_ap_vld(),
.ph_hit_o_0_12_6_V_ap_vld(),
.ph_hit_o_0_12_7_V_ap_vld(),
.ph_hit_o_0_12_8_V_ap_vld(),

// SHIFT LOGIC


// SHIFT LOGIC - INPUT: [time_i]

if (feed_in_time_i == 1'h1) begin
	for (i=0; i<7; i=i+1) begin
		for (j=0; j<9; j=j+1) begin
			for (k=0; k<2; k=k+1) begin
				if (k==0) begin
					if (j==0) begin
						if (i==0) begin
							reg_time_i[i][j][k] <= bus_time_i;
						end else begin
							reg_time_i[i][j][k] <= reg_time_i[i-1][9-1][2-1];
						end
					end else begin
						reg_time_i[i][j][k] <= reg_time_i[i][j-1][2-1];
					end
				end else begin
					reg_time_i[i][j][k] <= reg_time_i[i][j][k-1];
				end
			end
		end
	end
end else begin
	for (i=0; i<7; i=i+1) begin
		for (j=0; j<9; j=j+1) begin
			for (k=0; k<2; k=k+1) begin
				reg_time_i[i][j][k] <= reg_time_i[i][j][k];
			end
		end
	end
end

// SHIFT LOGIC - INPUT: [vl_i]

if (feed_in_vl_i == 1'h1) begin
	for (i=0; i<13; i=i+1) begin
		for (j=0; j<9; j=j+1) begin
			if (j==0) begin
				if (i==0) begin
					reg_vl_i[i][j] <= bus_vl_i;
				end else begin
					reg_vl_i[i][j] <= reg_vl_i[i-1][9-1];
				end
			end else begin
				reg_vl_i[i][j] <= reg_vl_i[i][j-1];
			end
		end
	end
end else begin
	for (i=0; i<13; i=i+1) begin
		for (j=0; j<9; j=j+1) begin
			reg_vl_i[i][j] <= reg_vl_i[i][j];
		end
	end
end

// SHIFT LOGIC - INPUT: [q_i]

if (feed_in_q_i == 1'h1) begin
	for (i=0; i<13; i=i+1) begin
		for (j=0; j<9; j=j+1) begin
			for (k=0; k<3; k=k+1) begin
				if (k==0) begin
					if (j==0) begin
						if (i==0) begin
							reg_q_i[i][j][k] <= bus_q_i;
						end else begin
							reg_q_i[i][j][k] <= reg_q_i[i-1][9-1][3-1];
						end
					end else begin
						reg_q_i[i][j][k] <= reg_q_i[i][j-1][3-1];
					end
				end else begin
					reg_q_i[i][j][k] <= reg_q_i[i][j][k-1];
				end
			end
		end
	end
end else begin
	for (i=0; i<13; i=i+1) begin
		for (j=0; j<9; j=j+1) begin
			for (k=0; k<3; k=k+1) begin
				reg_q_i[i][j][k] <= reg_q_i[i][j][k];
			end
		end
	end
end

// SHIFT LOGIC - INPUT: [cpatr_i]

if (feed_in_cpatr_i == 1'h1) begin
	for (i=0; i<6; i=i+1) begin
		for (j=0; j<9; j=j+1) begin
			for (k=0; k<2; k=k+1) begin
				if (k==0) begin
					if (j==0) begin
						if (i==0) begin
							reg_cpatr_i[i][j][k] <= bus_cpatr_i;
						end else begin
							reg_cpatr_i[i][j][k] <= reg_cpatr_i[i-1][9-1][2-1];
						end
					end else begin
						reg_cpatr_i[i][j][k] <= reg_cpatr_i[i][j-1][2-1];
					end
				end else begin
					reg_cpatr_i[i][j][k] <= reg_cpatr_i[i][j][k-1];
				end
			end
		end
	end
end else begin
	for (i=0; i<6; i=i+1) begin
		for (j=0; j<9; j=j+1) begin
			for (k=0; k<2; k=k+1) begin
				reg_cpatr_i[i][j][k] <= reg_cpatr_i[i][j][k];
			end
		end
	end
end

// SHIFT LOGIC - INPUT: [ph_i]

if (feed_in_ph_i == 1'h1) begin
	for (i=0; i<6; i=i+1) begin
		for (j=0; j<9; j=j+1) begin
			for (k=0; k<2; k=k+1) begin
				if (k==0) begin
					if (j==0) begin
						if (i==0) begin
							reg_ph_i[i][j][k] <= bus_ph_i;
						end else begin
							reg_ph_i[i][j][k] <= reg_ph_i[i-1][9-1][2-1];
						end
					end else begin
						reg_ph_i[i][j][k] <= reg_ph_i[i][j-1][2-1];
					end
				end else begin
					reg_ph_i[i][j][k] <= reg_ph_i[i][j][k-1];
				end
			end
		end
	end
end else begin
	for (i=0; i<6; i=i+1) begin
		for (j=0; j<9; j=j+1) begin
			for (k=0; k<2; k=k+1) begin
				reg_ph_i[i][j][k] <= reg_ph_i[i][j][k];
			end
		end
	end
end

// SHIFT LOGIC - INPUT: [th11_i]

if (feed_in_th11_i == 1'h1) begin
	for (i=0; i<6; i=i+1) begin
		for (j=0; j<9; j=j+1) begin
			for (k=0; k<2; k=k+1) begin
				if (k==0) begin
					if (j==0) begin
						if (i==0) begin
							reg_th11_i[i][j][k] <= bus_th11_i;
						end else begin
							reg_th11_i[i][j][k] <= reg_th11_i[i-1][9-1][2-1];
						end
					end else begin
						reg_th11_i[i][j][k] <= reg_th11_i[i][j-1][2-1];
					end
				end else begin
					reg_th11_i[i][j][k] <= reg_th11_i[i][j][k-1];
				end
			end
		end
	end
end else begin
	for (i=0; i<6; i=i+1) begin
		for (j=0; j<9; j=j+1) begin
			for (k=0; k<2; k=k+1) begin
				reg_th11_i[i][j][k] <= reg_th11_i[i][j][k];
			end
		end
	end
end

// SHIFT LOGIC - INPUT: [th_i]

if (feed_in_th_i == 1'h1) begin
	for (i=0; i<3; i=i+1) begin
		for (j=0; j<3; j=j+1) begin
			for (k=0; k<4; k=k+1) begin
				if (k==0) begin
					if (j==0) begin
						if (i==0) begin
							reg_th_i[i][j][k] <= bus_th_i;
						end else begin
							reg_th_i[i][j][k] <= reg_th_i[i-1][3-1][4-1];
						end
					end else begin
						reg_th_i[i][j][k] <= reg_th_i[i][j-1][4-1];
					end
				end else begin
					reg_th_i[i][j][k] <= reg_th_i[i][j][k-1];
				end
			end
		end
	end
end else begin
	for (i=0; i<3; i=i+1) begin
		for (j=0; j<3; j=j+1) begin
			for (k=0; k<4; k=k+1) begin
				reg_th_i[i][j][k] <= reg_th_i[i][j][k];
			end
		end
	end
end

// SHIFT LOGIC - INPUT: [phzvl_i]

if (feed_in_phzvl_i == 1'h1) begin
	for (i=0; i<13; i=i+1) begin
		for (j=0; j<9; j=j+1) begin
			if (j==0) begin
				if (i==0) begin
					reg_phzvl_i[i][j] <= bus_phzvl_i;
				end else begin
					reg_phzvl_i[i][j] <= reg_phzvl_i[i-1][9-1];
				end
			end else begin
				reg_phzvl_i[i][j] <= reg_phzvl_i[i][j-1];
			end
		end
	end
end else begin
	for (i=0; i<13; i=i+1) begin
		for (j=0; j<9; j=j+1) begin
			reg_phzvl_i[i][j] <= reg_phzvl_i[i][j];
		end
	end
end

// SHIFT LOGIC - INPUT: [ph_hit_i]

if (feed_in_ph_hit_i == 1'h1) begin
	for (i=0; i<13; i=i+1) begin
		for (j=0; j<9; j=j+1) begin
			if (j==0) begin
				if (i==0) begin
					reg_ph_hit_i[i][j] <= bus_ph_hit_i;
				end else begin
					reg_ph_hit_i[i][j] <= reg_ph_hit_i[i-1][9-1];
				end
			end else begin
				reg_ph_hit_i[i][j] <= reg_ph_hit_i[i][j-1];
			end
		end
	end
end else begin
	for (i=0; i<13; i=i+1) begin
		for (j=0; j<9; j=j+1) begin
			reg_ph_hit_i[i][j] <= reg_ph_hit_i[i][j];
		end
	end
end

// SHIFT LOGIC - OUTPUT: [time_o]

if (feed_out_time_o == 1'h1) begin
	for (i=0; i<1; i=i+1) begin
		for (j=0; j<7; j=j+1) begin
			for (k=0; k<9; k=k+1) begin
				for (l=0; l<2; l=l+1) begin
					if (l==0) begin
						if (k==0) begin
							if (j==0) begin
								if (i==0) begin
									reg_time_o[i][j][k][l] <= bus_time_o;
								end else begin
									reg_time_o[i][j][k][l] <= reg_time_o[i-1][7-1][9-1][2-1];
								end
							end else begin
								reg_time_o[i][j][k][l] <= reg_time_o[i][j-1][9-1][2-1];
							end
						end else begin
							reg_time_o[i][j][k][l] <= reg_time_o[i][j][k-1][2-1];
						end
					end else begin
						reg_time_o[i][j][k][l] <= reg_time_o[i][j][k][l-1];
						if (l==2-1 && k==9-1 && j==7-1 && i==1-1) begin
							bus_time_o <= reg_time_o[i][j][k][l];
						end
					end
				end
			end
		end
	end
end else if (load_out_time_o == 1'h1) begin
	for (i=0; i<1; i=i+1) begin
		for (j=0; j<7; j=j+1) begin
			for (k=0; k<9; k=k+1) begin
				for (l=0; l<2; l=l+1) begin
					reg_time_o[i][j][k][l] <= wire_time_o[i][j][k][l];
				end
			end
		end
	end
end else begin
	for (i=0; i<1; i=i+1) begin
		for (j=0; j<7; j=j+1) begin
			for (k=0; k<9; k=k+1) begin
				for (l=0; l<2; l=l+1) begin
					reg_time_o[i][j][k][l] <= reg_time_o[i][j][k][l];
				end
			end
		end
	end
	bus_time_o <= bus_time_o;
end

// SHIFT LOGIC - OUTPUT: [vl_o]

if (feed_out_vl_o == 1'h1) begin
	for (i=0; i<1; i=i+1) begin
		for (j=0; j<13; j=j+1) begin
			for (k=0; k<9; k=k+1) begin
				if (k==0) begin
					if (j==0) begin
						if (i==0) begin
							reg_vl_o[i][j][k] <= bus_vl_o;
						end else begin
							reg_vl_o[i][j][k] <= reg_vl_o[i-1][13-1][9-1];
						end
					end else begin
						reg_vl_o[i][j][k] <= reg_vl_o[i][j-1][9-1];
					end
				end else begin
					reg_vl_o[i][j][k] <= reg_vl_o[i][j][k-1];
					if (k==9-1 && j==13-1 && i==1-1) begin
						bus_vl_o <= reg_vl_o[i][j][k];
					end
				end
			end
		end
	end
end else if (load_out_vl_o == 1'h1) begin
	for (i=0; i<1; i=i+1) begin
		for (j=0; j<13; j=j+1) begin
			for (k=0; k<9; k=k+1) begin
				reg_vl_o[i][j][k] <= wire_vl_o[i][j][k];
			end
		end
	end
end else begin
	for (i=0; i<1; i=i+1) begin
		for (j=0; j<13; j=j+1) begin
			for (k=0; k<9; k=k+1) begin
				reg_vl_o[i][j][k] <= reg_vl_o[i][j][k];
			end
		end
	end
	bus_vl_o <= bus_vl_o;
end

// SHIFT LOGIC - OUTPUT: [q_o]

if (feed_out_q_o == 1'h1) begin
	for (i=0; i<1; i=i+1) begin
		for (j=0; j<13; j=j+1) begin
			for (k=0; k<9; k=k+1) begin
				for (l=0; l<3; l=l+1) begin
					if (l==0) begin
						if (k==0) begin
							if (j==0) begin
								if (i==0) begin
									reg_q_o[i][j][k][l] <= bus_q_o;
								end else begin
									reg_q_o[i][j][k][l] <= reg_q_o[i-1][13-1][9-1][3-1];
								end
							end else begin
								reg_q_o[i][j][k][l] <= reg_q_o[i][j-1][9-1][3-1];
							end
						end else begin
							reg_q_o[i][j][k][l] <= reg_q_o[i][j][k-1][3-1];
						end
					end else begin
						reg_q_o[i][j][k][l] <= reg_q_o[i][j][k][l-1];
						if (l==3-1 && k==9-1 && j==13-1 && i==1-1) begin
							bus_q_o <= reg_q_o[i][j][k][l];
						end
					end
				end
			end
		end
	end
end else if (load_out_q_o == 1'h1) begin
	for (i=0; i<1; i=i+1) begin
		for (j=0; j<13; j=j+1) begin
			for (k=0; k<9; k=k+1) begin
				for (l=0; l<3; l=l+1) begin
					reg_q_o[i][j][k][l] <= wire_q_o[i][j][k][l];
				end
			end
		end
	end
end else begin
	for (i=0; i<1; i=i+1) begin
		for (j=0; j<13; j=j+1) begin
			for (k=0; k<9; k=k+1) begin
				for (l=0; l<3; l=l+1) begin
					reg_q_o[i][j][k][l] <= reg_q_o[i][j][k][l];
				end
			end
		end
	end
	bus_q_o <= bus_q_o;
end

// SHIFT LOGIC - OUTPUT: [cpatr_o]

if (feed_out_cpatr_o == 1'h1) begin
	for (i=0; i<1; i=i+1) begin
		for (j=0; j<6; j=j+1) begin
			for (k=0; k<9; k=k+1) begin
				for (l=0; l<2; l=l+1) begin
					if (l==0) begin
						if (k==0) begin
							if (j==0) begin
								if (i==0) begin
									reg_cpatr_o[i][j][k][l] <= bus_cpatr_o;
								end else begin
									reg_cpatr_o[i][j][k][l] <= reg_cpatr_o[i-1][6-1][9-1][2-1];
								end
							end else begin
								reg_cpatr_o[i][j][k][l] <= reg_cpatr_o[i][j-1][9-1][2-1];
							end
						end else begin
							reg_cpatr_o[i][j][k][l] <= reg_cpatr_o[i][j][k-1][2-1];
						end
					end else begin
						reg_cpatr_o[i][j][k][l] <= reg_cpatr_o[i][j][k][l-1];
						if (l==2-1 && k==9-1 && j==6-1 && i==1-1) begin
							bus_cpatr_o <= reg_cpatr_o[i][j][k][l];
						end
					end
				end
			end
		end
	end
end else if (load_out_cpatr_o == 1'h1) begin
	for (i=0; i<1; i=i+1) begin
		for (j=0; j<6; j=j+1) begin
			for (k=0; k<9; k=k+1) begin
				for (l=0; l<2; l=l+1) begin
					reg_cpatr_o[i][j][k][l] <= wire_cpatr_o[i][j][k][l];
				end
			end
		end
	end
end else begin
	for (i=0; i<1; i=i+1) begin
		for (j=0; j<6; j=j+1) begin
			for (k=0; k<9; k=k+1) begin
				for (l=0; l<2; l=l+1) begin
					reg_cpatr_o[i][j][k][l] <= reg_cpatr_o[i][j][k][l];
				end
			end
		end
	end
	bus_cpatr_o <= bus_cpatr_o;
end

// SHIFT LOGIC - OUTPUT: [ph_o]

if (feed_out_ph_o == 1'h1) begin
	for (i=0; i<1; i=i+1) begin
		for (j=0; j<6; j=j+1) begin
			for (k=0; k<9; k=k+1) begin
				for (l=0; l<2; l=l+1) begin
					if (l==0) begin
						if (k==0) begin
							if (j==0) begin
								if (i==0) begin
									reg_ph_o[i][j][k][l] <= bus_ph_o;
								end else begin
									reg_ph_o[i][j][k][l] <= reg_ph_o[i-1][6-1][9-1][2-1];
								end
							end else begin
								reg_ph_o[i][j][k][l] <= reg_ph_o[i][j-1][9-1][2-1];
							end
						end else begin
							reg_ph_o[i][j][k][l] <= reg_ph_o[i][j][k-1][2-1];
						end
					end else begin
						reg_ph_o[i][j][k][l] <= reg_ph_o[i][j][k][l-1];
						if (l==2-1 && k==9-1 && j==6-1 && i==1-1) begin
							bus_ph_o <= reg_ph_o[i][j][k][l];
						end
					end
				end
			end
		end
	end
end else if (load_out_ph_o == 1'h1) begin
	for (i=0; i<1; i=i+1) begin
		for (j=0; j<6; j=j+1) begin
			for (k=0; k<9; k=k+1) begin
				for (l=0; l<2; l=l+1) begin
					reg_ph_o[i][j][k][l] <= wire_ph_o[i][j][k][l];
				end
			end
		end
	end
end else begin
	for (i=0; i<1; i=i+1) begin
		for (j=0; j<6; j=j+1) begin
			for (k=0; k<9; k=k+1) begin
				for (l=0; l<2; l=l+1) begin
					reg_ph_o[i][j][k][l] <= reg_ph_o[i][j][k][l];
				end
			end
		end
	end
	bus_ph_o <= bus_ph_o;
end

// SHIFT LOGIC - OUTPUT: [th11_o]

if (feed_out_th11_o == 1'h1) begin
	for (i=0; i<1; i=i+1) begin
		for (j=0; j<6; j=j+1) begin
			for (k=0; k<9; k=k+1) begin
				for (l=0; l<2; l=l+1) begin
					if (l==0) begin
						if (k==0) begin
							if (j==0) begin
								if (i==0) begin
									reg_th11_o[i][j][k][l] <= bus_th11_o;
								end else begin
									reg_th11_o[i][j][k][l] <= reg_th11_o[i-1][6-1][9-1][2-1];
								end
							end else begin
								reg_th11_o[i][j][k][l] <= reg_th11_o[i][j-1][9-1][2-1];
							end
						end else begin
							reg_th11_o[i][j][k][l] <= reg_th11_o[i][j][k-1][2-1];
						end
					end else begin
						reg_th11_o[i][j][k][l] <= reg_th11_o[i][j][k][l-1];
						if (l==2-1 && k==9-1 && j==6-1 && i==1-1) begin
							bus_th11_o <= reg_th11_o[i][j][k][l];
						end
					end
				end
			end
		end
	end
end else if (load_out_th11_o == 1'h1) begin
	for (i=0; i<1; i=i+1) begin
		for (j=0; j<6; j=j+1) begin
			for (k=0; k<9; k=k+1) begin
				for (l=0; l<2; l=l+1) begin
					reg_th11_o[i][j][k][l] <= wire_th11_o[i][j][k][l];
				end
			end
		end
	end
end else begin
	for (i=0; i<1; i=i+1) begin
		for (j=0; j<6; j=j+1) begin
			for (k=0; k<9; k=k+1) begin
				for (l=0; l<2; l=l+1) begin
					reg_th11_o[i][j][k][l] <= reg_th11_o[i][j][k][l];
				end
			end
		end
	end
	bus_th11_o <= bus_th11_o;
end

// SHIFT LOGIC - OUTPUT: [th_o]

if (feed_out_th_o == 1'h1) begin
	for (i=0; i<1; i=i+1) begin
		for (j=0; j<3; j=j+1) begin
			for (k=0; k<3; k=k+1) begin
				for (l=0; l<4; l=l+1) begin
					if (l==0) begin
						if (k==0) begin
							if (j==0) begin
								if (i==0) begin
									reg_th_o[i][j][k][l] <= bus_th_o;
								end else begin
									reg_th_o[i][j][k][l] <= reg_th_o[i-1][3-1][3-1][4-1];
								end
							end else begin
								reg_th_o[i][j][k][l] <= reg_th_o[i][j-1][3-1][4-1];
							end
						end else begin
							reg_th_o[i][j][k][l] <= reg_th_o[i][j][k-1][4-1];
						end
					end else begin
						reg_th_o[i][j][k][l] <= reg_th_o[i][j][k][l-1];
						if (l==4-1 && k==3-1 && j==3-1 && i==1-1) begin
							bus_th_o <= reg_th_o[i][j][k][l];
						end
					end
				end
			end
		end
	end
end else if (load_out_th_o == 1'h1) begin
	for (i=0; i<1; i=i+1) begin
		for (j=0; j<3; j=j+1) begin
			for (k=0; k<3; k=k+1) begin
				for (l=0; l<4; l=l+1) begin
					reg_th_o[i][j][k][l] <= wire_th_o[i][j][k][l];
				end
			end
		end
	end
end else begin
	for (i=0; i<1; i=i+1) begin
		for (j=0; j<3; j=j+1) begin
			for (k=0; k<3; k=k+1) begin
				for (l=0; l<4; l=l+1) begin
					reg_th_o[i][j][k][l] <= reg_th_o[i][j][k][l];
				end
			end
		end
	end
	bus_th_o <= bus_th_o;
end

// SHIFT LOGIC - OUTPUT: [phzvl_o]

if (feed_out_phzvl_o == 1'h1) begin
	for (i=0; i<1; i=i+1) begin
		for (j=0; j<13; j=j+1) begin
			for (k=0; k<9; k=k+1) begin
				if (k==0) begin
					if (j==0) begin
						if (i==0) begin
							reg_phzvl_o[i][j][k] <= bus_phzvl_o;
						end else begin
							reg_phzvl_o[i][j][k] <= reg_phzvl_o[i-1][13-1][9-1];
						end
					end else begin
						reg_phzvl_o[i][j][k] <= reg_phzvl_o[i][j-1][9-1];
					end
				end else begin
					reg_phzvl_o[i][j][k] <= reg_phzvl_o[i][j][k-1];
					if (k==9-1 && j==13-1 && i==1-1) begin
						bus_phzvl_o <= reg_phzvl_o[i][j][k];
					end
				end
			end
		end
	end
end else if (load_out_phzvl_o == 1'h1) begin
	for (i=0; i<1; i=i+1) begin
		for (j=0; j<13; j=j+1) begin
			for (k=0; k<9; k=k+1) begin
				reg_phzvl_o[i][j][k] <= wire_phzvl_o[i][j][k];
			end
		end
	end
end else begin
	for (i=0; i<1; i=i+1) begin
		for (j=0; j<13; j=j+1) begin
			for (k=0; k<9; k=k+1) begin
				reg_phzvl_o[i][j][k] <= reg_phzvl_o[i][j][k];
			end
		end
	end
	bus_phzvl_o <= bus_phzvl_o;
end

// SHIFT LOGIC - OUTPUT: [ph_hit_o]

if (feed_out_ph_hit_o == 1'h1) begin
	for (i=0; i<1; i=i+1) begin
		for (j=0; j<13; j=j+1) begin
			for (k=0; k<9; k=k+1) begin
				if (k==0) begin
					if (j==0) begin
						if (i==0) begin
							reg_ph_hit_o[i][j][k] <= bus_ph_hit_o;
						end else begin
							reg_ph_hit_o[i][j][k] <= reg_ph_hit_o[i-1][13-1][9-1];
						end
					end else begin
						reg_ph_hit_o[i][j][k] <= reg_ph_hit_o[i][j-1][9-1];
					end
				end else begin
					reg_ph_hit_o[i][j][k] <= reg_ph_hit_o[i][j][k-1];
					if (k==9-1 && j==13-1 && i==1-1) begin
						bus_ph_hit_o <= reg_ph_hit_o[i][j][k];
					end
				end
			end
		end
	end
end else if (load_out_ph_hit_o == 1'h1) begin
	for (i=0; i<1; i=i+1) begin
		for (j=0; j<13; j=j+1) begin
			for (k=0; k<9; k=k+1) begin
				reg_ph_hit_o[i][j][k] <= wire_ph_hit_o[i][j][k];
			end
		end
	end
end else begin
	for (i=0; i<1; i=i+1) begin
		for (j=0; j<13; j=j+1) begin
			for (k=0; k<9; k=k+1) begin
				reg_ph_hit_o[i][j][k] <= reg_ph_hit_o[i][j][k];
			end
		end
	end
	bus_ph_hit_o <= bus_ph_hit_o;
end

// RESET LOGIC

for (i=0; i<7; i=i+1) begin
	for (j=0; j<9; j=j+1) begin
		for (k=0; k<2; k=k+1) begin
			reg_time_i[i][j][k] <= 0;
		end
	end
end
for (i=0; i<13; i=i+1) begin
	for (j=0; j<9; j=j+1) begin
		reg_vl_i[i][j] <= 0;
	end
end
for (i=0; i<13; i=i+1) begin
	for (j=0; j<9; j=j+1) begin
		for (k=0; k<3; k=k+1) begin
			reg_q_i[i][j][k] <= 0;
		end
	end
end
for (i=0; i<6; i=i+1) begin
	for (j=0; j<9; j=j+1) begin
		for (k=0; k<2; k=k+1) begin
			reg_cpatr_i[i][j][k] <= 0;
		end
	end
end
for (i=0; i<6; i=i+1) begin
	for (j=0; j<9; j=j+1) begin
		for (k=0; k<2; k=k+1) begin
			reg_ph_i[i][j][k] <= 0;
		end
	end
end
for (i=0; i<6; i=i+1) begin
	for (j=0; j<9; j=j+1) begin
		for (k=0; k<2; k=k+1) begin
			reg_th11_i[i][j][k] <= 0;
		end
	end
end
for (i=0; i<3; i=i+1) begin
	for (j=0; j<3; j=j+1) begin
		for (k=0; k<4; k=k+1) begin
			reg_th_i[i][j][k] <= 0;
		end
	end
end
for (i=0; i<13; i=i+1) begin
	for (j=0; j<9; j=j+1) begin
		reg_phzvl_i[i][j] <= 0;
	end
end
for (i=0; i<13; i=i+1) begin
	for (j=0; j<9; j=j+1) begin
		reg_ph_hit_i[i][j] <= 0;
	end
end
for (i=0; i<1; i=i+1) begin
	for (j=0; j<7; j=j+1) begin
		for (k=0; k<9; k=k+1) begin
			for (l=0; l<2; l=l+1) begin
				reg_time_o[i][j][k][l] <= 0;
			end
		end
	end
end
bus_time_o <= 0;
for (i=0; i<1; i=i+1) begin
	for (j=0; j<13; j=j+1) begin
		for (k=0; k<9; k=k+1) begin
			reg_vl_o[i][j][k] <= 0;
		end
	end
end
bus_vl_o <= 0;
for (i=0; i<1; i=i+1) begin
	for (j=0; j<13; j=j+1) begin
		for (k=0; k<9; k=k+1) begin
			for (l=0; l<3; l=l+1) begin
				reg_q_o[i][j][k][l] <= 0;
			end
		end
	end
end
bus_q_o <= 0;
for (i=0; i<1; i=i+1) begin
	for (j=0; j<6; j=j+1) begin
		for (k=0; k<9; k=k+1) begin
			for (l=0; l<2; l=l+1) begin
				reg_cpatr_o[i][j][k][l] <= 0;
			end
		end
	end
end
bus_cpatr_o <= 0;
for (i=0; i<1; i=i+1) begin
	for (j=0; j<6; j=j+1) begin
		for (k=0; k<9; k=k+1) begin
			for (l=0; l<2; l=l+1) begin
				reg_ph_o[i][j][k][l] <= 0;
			end
		end
	end
end
bus_ph_o <= 0;
for (i=0; i<1; i=i+1) begin
	for (j=0; j<6; j=j+1) begin
		for (k=0; k<9; k=k+1) begin
			for (l=0; l<2; l=l+1) begin
				reg_th11_o[i][j][k][l] <= 0;
			end
		end
	end
end
bus_th11_o <= 0;
for (i=0; i<1; i=i+1) begin
	for (j=0; j<3; j=j+1) begin
		for (k=0; k<3; k=k+1) begin
			for (l=0; l<4; l=l+1) begin
				reg_th_o[i][j][k][l] <= 0;
			end
		end
	end
end
bus_th_o <= 0;
for (i=0; i<1; i=i+1) begin
	for (j=0; j<13; j=j+1) begin
		for (k=0; k<9; k=k+1) begin
			reg_phzvl_o[i][j][k] <= 0;
		end
	end
end
bus_phzvl_o <= 0;
for (i=0; i<1; i=i+1) begin
	for (j=0; j<13; j=j+1) begin
		for (k=0; k<9; k=k+1) begin
			reg_ph_hit_o[i][j][k] <= 0;
		end
	end
end
bus_ph_hit_o <= 0;
